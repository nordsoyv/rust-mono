title "copy of 231 II"

// workaround to avoid Compiler Error for config access block
config pulse

config hub {
  hub: 14900
  table accounts = custom.Account_2      //accounts custom table
  table survey = p1850259384.response  //relationship survey
  table contacts = p1862934241.response
  table healthCheck = p1860215844.response      //healthcheck survey
  table cases = am.CASE
  table respondent = p1850259384.respondent
  table revenue = custom.Historical_Revenue  // historical revenue custom table.
  table new = custom.Account_2
  table ejournal = custom.eJournal


// config report cr {
//   currentPeriod: InMonth(survey:interview_start,-1,0)
//   previousPeriod: InMonth(survey:interview_start,-13,-11)
//    // <-- unmatching brackets in comments

  //accounts --> revenue
  relation oneToMany #rel3 {
    primaryKey: accounts:accountID
    foreignKey: revenue:accountID
  }

  // accounts --> Health
  relation oneToMany #rel2 {
    primaryKey: accounts:AccountID
    foreignKey: healthCheck:shortAccountID

  }
  // accounts --> contact db --> survey
  relation oneToMany #rel4 {
    primaryKey: accounts:AccountID
    foreignKey: contacts:shortAccountID
  }
  //accounts --> eJournal
  relation oneToMany #rel5 {
    primaryKey: accounts:eJournalAccountNumber
    foreignKey: ejournal:compid
  }

}
layoutArea toolbar {
  filter multiselect #accountOwenr {
    label: "Account Owner"
    optionsFrom: accounts:AccountOwner
  }
  filter multiselect #risk {
    label: "Revenue Risk"
    filterType: postAggregate
    option checkbox #a {
      label: "High"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10
    }
    option checkbox #b {
      label: "Medium"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(respondent:respid) * 100 > 4 AND average(SCORE(survey:Q1)) < 7 OR average(SCORE(healthCheck:NPS)) < 5
    }
    option checkbox #c {
      label: "Low"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(respondent:respid) * 100 > 4 AND average(SCORE(survey:Q1)) > 6 AND count(healthCheck:responseid) > 0 AND average(SCORE(healthCheck:NPS)) > 6 OR count(healthCheck:responseid) > 0
    }
  }

  filter multiselect #region {
    label: "Region"
    optionsFrom: accounts:SalesRegion
  }

  filter multiselect #role {
    label: "Role"
    option checkbox #r1 {
      label: "Decision maker"
      value: contacts:contactRole = "Decision maker"
    }
    option checkbox #r2 {
      label: "Influencer"
      value: contacts:contactRole = "Influencer"
    }

  }
  filter multiselect #period {
    label: "Reporting period"
    option checkbox #s1 {
      label: "Last quarter"
      value: survey:interview_start > 2017-09-30 AND survey:interview_start < 2018-01-01
    }
    option checkbox #s2 {
      label: "Last 6 months"
      value: survey:interview_start > 2017-10-23
    }
    option checkbox #s3 {
      label: "Last 12 months"
      value: survey:interview_start > 2017-01-23
    }
  }

  filter multiselect #renewal {
    label: "Renewal period"
    option checkbox #q1 {
      label: "Q1 2018"
      value: accounts:RenewalDate > 2018-01-01 AND accounts:RenewalDate < 2018-04-01
    }
    option checkbox #q2 {
      label: "Q2 2018"
      value: accounts:RenewalDate > 2018-03-31 AND accounts:RenewalDate < 2018-07-01
    }
    option checkbox #q3 {
      label: "Q3 2018"
      value: accounts:RenewalDate > 2018-06-30 AND accounts:RenewalDate < 2018-10-01
    }
    option checkbox #q4 {
      label: "Q4 2018"
      value: accounts:RenewalDate > 2018-09-30 AND accounts:RenewalDate < 2019-01-01
    }
  }
}

custom properties #cp {
  // variables to be used by writing e.g. @cp.revenueRiskValue // cr =
  revenueRiskValue: IIF((sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10, 3, IIF((sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < 10, 2, 1))
}

config report #cr {
  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Confirmit%20Demo/confirmit3Dlogo.jpg"
  formatter date #date11 {
    shortForm: true
    emptyValue: "None"
  }
  formatter date #dateFormat {
    inputFormat: "YYYYMM"
    formatString: "MMM"
  }
  formatter date #date12 {
    locale: en
    //format: "DD MMMM YYYY"
    shortForm: false
  }
  formatter value #valueFMT {
    emptyValue: " "
  }
  formatter number #formatterID {
    numberDecimals: 0
    prefix: "$ "
    decimalSeparator: "."
    integerSeparator: " "
    shortForm: true
  }
  formatter number #formatterLTR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    emptyValue: "-"
  }
  formatter number #formatterRR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    postfix: " %"
  }

  formatter color #formatterColor {
    thresholds: #009900 >=9 , #b34700 >=7, #b30000 >=0
  }
  formatter color #formatterColor2 {
    thresholds: #0099AA >=9 , #b347AA >=7, #b300AA >=0
  }
  formatter number #metricFormat {
    numberDecimals: 1
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
  }

  formatter number #responsesFormat {
    numberDecimals: 0
    shortForm: false
  }
  // duplicate
  // formatter date dateFormat {
  //   inputFormat: "YYYYMM"
  //   formatString: "MMM YY"
  // }

  formatter color #riskStringFormatter {
    thresholds: Unknown = 0 , Low = 1, Medium = 2, High = 3
  }

  formatter color #riskBgColorFormatter {
    thresholds: #23C813 >= 9, #FFAB00 >= 7, #ff0000 >= 0
  }
  formatter color #risk {
    thresholds: #23C813 >= 9, #FFAB00 >= 7, #ff0000 >= 0
  }

  formatter color #backgroundColor {
    thresholds: #e8f8e0 >= 9, #ffeed6 >= 7, #fedfe2 >= 0
  }
  formatter color #valueColor {
    thresholds: #388e3c >= 9, #ff6d00 >= 7, #d40000 >= 0
  }
  formatter color #valueColorFormatter {
    thresholds: #5ba35d >= 8.5, #ffa156 >= 6.5, #dd3435 >= 0
  }
  formatter objectProperty #textPicker {
    property: text
  }

  formatter color #riskColorFormatter {
    thresholds: #FA5263 >= 99%, #FFBD5B >=49%, #82D854 >0%
  }
  ltrTarget: 9

  view metric #metrics {
    valueColorFormatter: valueColor
    fontSize: large
    backgroundColorFormatter: transparent
  }
  view metricWithChange #metricsWithChange {
    backgroundColorFormatter: backgroundColor
    valueColorFormatter: valueColor
    fontSize: small
    roundCorners: true
  }
}

page #Overview {
  label: "Overview"

  widget kpi {
    label: "Global NPS"
    size: small
    tile kpi {
      label: "NPS"
      value: NPS(survey:Q1) * 100
      min: -100
      max: 100
      format: formatterLTR
      targetFormat: formatterLTR
      gaugeColorFormat: riskBgColorFormatter  // valueColor
      tile value {
        label: "Responses"
        value: count(survey:Q1)
        max: count(survey:responseid)
        format: integer
      }
      tile value {
        label: "Yearly change"
        //value: average(score(survey:Q1),@cr.currentPeriodFilter)-average(score(survey:Q1),@cr.previousPeriodFilter)
        format: formatterLTR
      }
    }
  }
  widget portfolioBreakdown {
    label: "Average LTR monthly"
    size: small

    category: calendarMonth(survey:interview_start)
    categoryFormat: dateFormat
    value: average(score(survey:Q1))
    format: formatterLTR
  }
  widget kpi {
    label: "Overall Satisfaction"
    size: small
    tile kpi {
      label: "AVG"
      value: average(score(survey:Q1))
      min: 0
      max: 10
      format: formatterLTR
      targetFormat: formatterLTR
      gaugeColorFormat: kpiColorFormatter       //valueColor
      tile value {
        label: "Responses"
        value: count(survey:responseid, survey:status = "Complete")// AND @cp.currentPeriodFilter)
        max: count(survey:responseid)
        format: integer
      }
      tile value {
        label: "Yearly change"
        value: average(score(survey:Q4)) - average(score(survey:Q4))
        format: formatterLTR
      }
    }
  }

  widget kpi {
    label: "Internal View"
    size: small
    tile kpi {
      label: "AVG"
      value: average(score(healthCheck:Q1))
      min: 0
      max: 10
      format: formatterLTR
      targetFormat: formatterLTR
      gaugeColorFormat: kpiColorFormatter       //valueColor
    }
  }

  widget portfolioBreakdown #R {
    label: "Portfolio Risk Assessment"
    size: medium
    category: CalendarMONTH(accounts:RenewalDate)
    segment: IIF(count(healthCheck:responseid, true, accounts:) > 0, IIF(average(SCORE(healthCheck:Q2), true, accounts:) >= 9, "Medium", IIF(average(SCORE(healthCheck:Q2), true, accounts:) >= 5, "High", "Unknown")), "Safe")
    value: count(survey:responseid)
  }

  widget markdown {
    size: small

    markdown: "
## Churn Risk assessment model
The Risk is calculated from the NPS score and Internal Account Check score
The following Risk model is applied
A score between 0 and 6 indicates High risk of churn
A score between 7 and 8 indicates Medium risk
A score between 9 and 10 indicate that account is Safe.

in case of lacking responses the risk is unknown"
  }

  widget recentResponses #yy {
    label: "Customer Responses"
    showHeader: true
    view comment #fff {
      lines: 3
    }
    size: medium
    table: survey:
    view metric #metrics {
      valueColorFormatter: valueColor
      fontSize: large
      backgroundColorFormatter: transparent
    }
    column response #x1 {
      sortBy: footer
      footer: survey:interview_end
      header: survey:FirstName + " " + survey:LastName + " - " + accounts:AccountName
      comment: survey:Q2
      commentFormat: commentFormat
      navigateTo: Contact
    }
    column metric #ltr2 {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      target: 10
      view: metrics
    }
  }
  widget recentResponses #IV {
    label: "Internal View Responses"
    table: healthCheck:
    size: small
    lines: 3
    view metric #metrics {
      valueColorFormatter: valueColor
      fontSize: large
      backgroundColorFormatter: transparent
    }
    column response {
      sortBy: footer
      footer: healthCheck:interview_end
      header: AnswerText(accounts:AccountOwner) + " - " + AnswerText(accounts:SalesRegion)
      comment: healthCheck:Q3

    }
    column metric #ltr3 {
      label: "LTR  Estimate"
      value: average(score(healthCheck:Q2))
      target: 9
      view: metrics
    }
  }

  widget topAccounts {
    table: accounts:
    size: small
    sortColumn: main
    navigateTo: Account
    hierarchy: accounts:ParentAccountID
    view metricWithChange #metrics {
      valueColorFormatter: valueColor
      backgroundColorFormatter: transparent
      fontSize: medium
    }
    column accounts #main {
      accountName: accounts:AccountName
      revenue: SUM(accounts:AnnualAccountValue)
      value: SUM(accounts:AnnualAccountValue)
    }
    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      // previous: average(score(survey:Q1))
      //value: average(score(survey:Q1) @cr.currentPeriodFilter)
      // previous: average(score(survey:Q1),@cr.previousPeriodFilter)
      format: formatterLTR
      target: @cr.ltrTarget
      view: metrics
    }
  }
  widget portfolioBreakdown {
    label: "NPS Breakdown by Role (%)"
    size: medium

    category: contacts:ContactRole
    segment: survey:NPSSegment
    value: count(survey:responseId)

    percent: on
    // palette: @cp.palette
    // format: floatNumber
  }

  widget portfolioBreakdown {
    label: "NPS Breakdown by Role"
    size: medium

    category: contacts:ContactRole
    segment: survey:NPSSegment
    value: count(survey:responseId)

    percent: off
  }
}

page #AccountRiskFactors {
  label: "Account Risk Factors"

  widget markdown {
    size: medium

    markdown: "
## Confirmit Confidential Information
Please do not use this report in the external demos"
  }
  widget accountList {
    label: "Accounts"
    table: accounts:
    sortColumn: accountName
    //sortOrder: accending
    navigateTo: Account
    size: large

    hierarchy: accounts:ParentAccountID

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
      //roundCorners:true
    }

    column hierarchy #accountName {
      label: "Account Name "
      value: accounts:AccountName
      rowHeader: true
    }

    column metric #ltr {
      label: "Client View"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column metric #hh {
      label: "Internal View"
      value: average(score(healthCheck:Q2))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column value #accountMan {
      label: "Account Owner"
      value: accounts:AccountOwner
    }

    column value #revRisk {
      label: "Revenue Risk " //Churn Risk
      value: @cp.revenueRiskValue
      align: center
      format: riskStringFormatter
    }
    column value #rev2017 {
      label: "2017 rev"
      value: sum(revenue:AnnualRevenue, revenue:year = 2017)
      format: formatterID
      align: right
    }
    column value #rev2016 {
      label: "2016 rev"
      value: sum(revenue:AnnualRevenue, revenue:year = 2016)
      format: formatterID
      align: right
    }
    column value #revDiff {
      label: "Rev diff"
      value: sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)
      format: formatterID
      align: right
    }
    column value #revDiffPercentage {
      label: "Rev diff"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100
      format: formatterRR
      align: right
    }
    column value #tickets {
      label: "eJournal total"
      value: sum(ejournal:closedTickets)
    }
    column value #ticketsOpen {
      label: "eJournal Open"
      value: sum(ejournal:openTickets)
    }

    column value #case2 {
      label: "Cases"
      value: COUNT(cases:CaseId)
      align: center
      format: responsesFormat

    }
    column value #responses {
      label: "Responses "
      format: valueFMTnses
      value: COUNT(survey:responseid, survey:status = "complete") //OR survey:status="incomplete"
      align: center
    }

    column value #rate {
      label: "Response Rate"
      value: COUNT(survey:responseId, survey:status = "complete" OR survey:status = "incomplete") * 100 / COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
      format: formatterRR
      align: center
    }
    column value #noResp {
      label: "No Response"
      value: COUNT(respondent:respid, respondent:smtpstatus = "messagesent") - COUNT(survey:responseid, survey:status = "Complete")
      align: center
    }
  }
}

page account #Account {
  label: "Account"


  widget search {
    table: accounts:
    layoutArea: "header"
    value: accounts:AccountName + " " + accounts:AccountId
    navigateTo: AccountPage
    iconType: "account"
  }


  widget title {
    table: accounts:
    layout column {
      tile value #c {
        value: accounts:accountName
      }
    }
  }

  widget summary {
    size: large
    table: accounts:

    tile metric {
      label: "LTR Average"
      value: average(score(survey:Q1))
      target: 7
    }

    tile metric {
      label: "Health check"
      value: average(score(healthCheck:Q2))
      target: 5
    }


    tile risk {
      label: "Revenue Risk"
        // need to tune formatting! add calculation
      value: @cp.revenueRiskValue
      textValue: IIF(@cp.revenueRiskValue = 3, "High", IIF(@cp.revenueRiskValue = 2, "Medium", IIF(@cp.revenueRiskValue = 1, "Low", "Unknown")))
      min: 1
      max: 3
      target: 0
      renewal: accounts:RenewalDate
      revenue: sum(revenue:AnnualRevenue, revenue:year = 2017)
      backgroundColorFormatter: riskColorFormatter
    }

    tile responseRate {
      invites: COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
      responses: COUNT(survey:responseId, survey:status = "complete" OR survey:status = "incomplete")
    }

    tile casesStatus {
      label: "Cases"
      open: COUNT(cases:CaseId)
      overdue: 0
    }
  }

  widget contactList #hg {
    size: large
    label: "Contacts "
    table: contacts:
    sortColumn: name
    sortOrder: descending
    navigateTo: Contact

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    view metric #ccc {
      valueColorFormatter: valueCases
    }
    column value #name {
      label: "Name"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #company {
      label: "Company"
      value: contacts:AccountName
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }

    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
    }
    column value #openCases {
      label: "Cases"
      value: COUNT(cases:CaseId)
      view: ccc
    }
    column value #lastResponse {
      label: "Last response "
      value: LAST(survey:interview_start, survey:interview_start)
      format: date11
      asign: center
    }
    column value #comments {
      label: "Comments"
      value: LAST(survey:Q2, survey:interview_start)
    }
  }

  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Date"
      value: cases:DateCreated
      align: center
      format: date12
    }

    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000818", "Health Check : At Risk", IIF(cases:Workflow = "1000819", "Health Check : High Potential", "Relationship : Recommend and/or Tech Detractors")))
    }
    column value #res {
      label: "Resolution"
      value: IIF(cases:lk_1548 = "5218" OR cases:lk_1548 = "5219" OR cases:lk_1548 = "5220", "Client specific", IIF(cases:lk_1548 = "5221" OR cases:lk_1548 = "5222" OR cases:lk_1548 = "5223", "Generic", IIF(cases:lk_1548 = "8319" OR cases:lk_1548 = "8320" OR cases:lk_1548 = "8321" OR cases:lk_1548 = "8322", "At risk: Action Taken", IIF(cases:lk_1548 = "8323" OR cases:lk_1548 = "8324", "High potential", "To Be Coded"))))
    }

    column value #link {

      label: "Action"
      value: cases:CaseLink
      view: link1
    }

  }
}

page contact #Contact {
  label: "Contact"


  widget search {
    table: contacts:
    layoutArea: "header"
    value: contacts:client_first_name + " " + contacts:client_last_name
    navigateTo: ContactList
  }



  widget title {
    view icon #icon {
      size: "60"
      roundedCorner: true
    }
    table: contacts:
    layout column {
      tile icon {
        value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/magdalenas/defaultLogo.PNG"//"http://is1.mzstatic.com/image/thumb/Purple71/v4/89/51/f4/8951f4f1-fd6b-fa59-38b2-191140473b9a/source/175x175bb.jpg"
      }
    }
    layout column {
      layout row {
        tile value {
          value: contacts:FirstName + " " + contacts:LastName
        }
        tile role {
          value: contacts:ContactRole
        }
      }
      layout row {
        tile company {
          value: contacts:AccountName
        }
      }
    }
  }

  widget summary {
    size: large
    table: contacts:
    tile contactDetails #cc {
      title: contacts:Title
      role: contacts:ContactRole
      email: contacts:email
      phone: contacts:Phone
      industry: contacts:Industry
    }

    tile accountDetails #cc4 {
      accountOwner: contacts:AccountOwner
      salesManager: contacts:SalesLeader1
      region: contacts:WorldRegion
      revenue: contacts:AnnualAccountValue
      renewalDate: accounts:RenewalDate

    }

    tile metric #a {
      label: "LTR"
      value: average(score(survey:Q1))
      target: 9
    }

    tile metric #da {
      label: "Surveys"
      value: count(survey:responseid)
    }

    tile casesStatus {
      label: Cases
      open: count(cases:CaseId)
      overdue: 0
    }
  }

  widget contactSurveys {
    label: "Surveys"
    table: survey:
    sortColumn: surveyDate
    sortOrder: ascending
    size: large
    navigateTo: SurveyResponse

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
      //roundCorners:true
    }

    column value #status {
      label: "Status"
      value: survey:status
      format: textPicker
    }


    column date #surveyDate {
      label: "Date"
      value: survey:interview_end

    }

    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column value #case2 {
      label: "Cases"
      value: COUNT(cases:CaseId)
      align: center
      format: responsesFormat
    }

    column value #comments {
      label: "Comments"
      value: survey:Q2
    }
  }

  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending
    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Date"
      value: cases:DateCreated
      align: center
      format: date12
    }

    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000818", "Health Check : At Risk", IIF(cases:Workflow = "1000819", "Health Check : High Potential", "Relationship : Recommend and/or Tech Detractors")))
    }
    column value #res {
      label: "Resolution"
      value: IIF(cases:lk_1548 = "5218" OR cases:lk_1548 = "5219" OR cases:lk_1548 = "5220", "Client specific", IIF(cases:lk_1548 = "5221" OR cases:lk_1548 = "5222" OR cases:lk_1548 = "5223", "Generic", IIF(cases:lk_1548 = "8319" OR cases:lk_1548 = "8320" OR cases:lk_1548 = "8321" OR cases:lk_1548 = "8322", "At risk: Action Taken", IIF(cases:lk_1548 = "8323" OR cases:lk_1548 = "8324", "High potential", "To Be Coded"))))
    }

    column value #link {

      label: "CaseLink"
      value: cases:CaseLink
      view: link1
    }
    widget contactSurveys {
      label: "Surveys"
      table: survey:
      sortColumn: is
      size: large
      navigateTo: SurveyResponse
      sortOrder: ascending
      view metricWithChange #metrics {
        backgroundColorFormatter: backgroundColor
        valueColorFormatter: valueColor
        fontSize: small
        roundCorners: true
      }
      column value {
        label: "Survey"
        value: "Relationship Survey"
      }
      column value #s2 {
        label: "Status"
        value: survey:status
      }
      column value #is {
        label: "Date"
        value: survey:interview_start
        format: dateRelative
      }
      column metric #s3 {
        label: "LTR"
      // value: average(score(survey:Q1), @cr.currentPeriodFilter)
      // previous: average(score(survey:Q1), @cr.previousPeriodFilter)
        target: @cr.ltrTarget
        format: formatterLTR
        align: center
        view: metrics
      }

      column value #s6 {
        label: "Comments"
        value: Last(survey:Q8, survey:interview_end)
      }
      view link #viewResp {
        label: "View Response"
      }
      column value {
        label: "Actions"
        value: 1
        view: viewResp
      }
    }

  }
  page #SurveyResponse {
    widget contactSurveyResponse {
      view title #defaultSurveyResponseTitle {
      }


      size: medium
      surveyResponseTitle {
        contactName: contacts:FirstName + " " + contacts:LastName
        surveyName: survey:SurveyId
        tile title #rt {
          contactName: contacts:FirstName + " " + contacts:LastName
          surveyName: survey:responseid
          view: defaultSurveyResponseTitle
        }
      }
      summary {
        rows: 4

        tile list #list1 {
          item value {
            value: survey:UploadedDate
            label: "Received"
            format: DDMMMYYYY
          }
          item value {
            value: survey:status
            label: "Status"
          }
          item email {
            value: survey:interview_start
            label: "Interview Start"
          }
          item value {
            value: survey:interview_end
            label: "Interview End"
          }
        }
        tile list #list2 {
          item value {
            value: "Relationship Survey"
            label: "Source"
          }
          item email {
            value: survey:responseid
            label: "Response ID"
          }
          item value {
            value: contacts:contactid
            label: "Respondent ID"
          }
        }
      }

      tab {
        label: "All"
        tile list {
          label: " "
          item comment {
            label: "First Name"
            value: accounts:FirstName
          }
          item comment {
            label: "Last Name"
            value: contacts:LastName
          }
          item comment {
            label: "Company name"
            value: accounts:AccountName
          }
          item comment {
            label: "Title"
            value: contacts:Title
          }
          item comment {
            label: "Role"
            value: contacts:ContactRole
          }
          view: defaulViewForListTile
        }
        tile list {
          label: "Key Metrics"
          item bar {
            label: "Likelihood to Recommend"
            value: average(score(survey:Q1))
          }
          item bar {
            label: "Overall Satisfaction"
            value: average(score(survey:Q4))
          }
          item comment {
            label: "Satisfaction with Technology"
            value: survey:Q8
          }
          view: defaulViewForListTile
        }
        tile list {
          label: "Product Satisfaction"
          item bar {
            label: "Technology"
            value: average(score(survey:Q7))
          }
          item bar {
            label: "Product is scalable"
            value: average(score(survey:Q9.1))
          }
          item bar {
            label: "Product is easy to use"
            value: average(score(survey:Q9.2))
          }
          item bar {
            label: "Product delivers results"
            value: average(score(survey:Q9.3))
          }
          view: defaulViewForListTile
        }
        tile list {
          label: "Service Satisfaction"
          item bar {
            label: "Provide Added Value"
            value: average(score(survey:Q3))
          }
          item bar {
            label: "Support business needs"
            value: average(score(survey:Q12))
          }
          view: defaulViewForListTile
        }
      }
      tab {
        label: "Comments"
        tile list {
          label: "Key"
          item comment {
            label: "label1"
            value: survey:Q2
          }
          item comment {
            label: "label2"
            value: survey:Q6
          }
        }
        view: defaulViewForListTile
      }
      tab {
        label: "CASE DATA"
        tile list {
          label: "NPS Detractor Alert"
          item bar {
            label: "Likelyhood to Recommend"
            value: average(score(survey:Q1))
          }
          item bar {
            label: "Overall Satisfaction"
            value: average(score(survey:Q4))
          }
          item comment {
            label: "Satisfaction with Technology"
            value: survey:Q8
          }
          view: defaulViewForListTile
        }
        tile list {
          label: "Product Satisfaction"
          item bar {
            label: "Technology"
            value: average(score(survey:Q7))
          }
          item bar {
            label: "Product is scalable"
            value: average(score(survey:Q9.1))
          }
          item bar {
            label: "Product is easy to use"
            value: average(score(survey:Q9.2))
          }
          item bar {
            label: "Product delivers results"
            value: average(score(survey:Q9.3))
          }
          view: defaulViewForListTile
        }
        tile list {
          label: "Service Satisfaction"
          item bar {
            label: "Provide Added Value"
            value: average(score(survey:Q3))
          }
          item bar {
            label: "Support business needs"
            value: average(score(survey:Q12))
          }
          view: defaulViewForListTile
        }
      }
    }
  }
}

title "VOC mch test"
config hub {
  hub: 14900
  table accounts = custom.Account_2
  table survey = p1850259384.response
  table surveyR = p1850259384.respondent
  table contacts = p1862934241.response
  table healthCheck = p1860215844.response      //healthcheck survey
  table health = p1860215844.response
  table cases = am.CASE
  table revenue = custom.Historical_Revenue
  table ejournal = custom.eJournal
  relation oneToMany #rel3 {
    primaryKey: accounts:accountID
    foreignKey: revenue:accountID
  }
  relation oneToMany #rel2 {
    primaryKey: accounts:AccountID
    foreignKey: healthCheck:shortAccountID
  }
  relation oneToMany #rel4 {
    primaryKey: accounts:AccountID
    foreignKey: contacts:shortAccountID
  }
  relation oneToMany #rel5 {
    primaryKey: accounts:eJournalAccountNumber
    foreignKey: ejournal:compid
  }

  variable auto #NAcc {
    label: "Real"
    table: accounts:
    value: accounts:TotalAccountValue
  }
  variable auto #NN {
    table: accounts:
    value: COUNT(survey:)
  }
  variable singleChoice #oo {
    label: "oo"
    table: accounts:
    option code {
      code: "Safe"
      score: 1
      label: "Safe"
    }
    option code {
      code: "Medium"
      score: 2
      label: "Medium"
    }
    option code {
      code: "High"
      score: 3
      label: "High"
    }
    option code {
      code: "Unknown"
      score: 4
      label: "Unknown"
    }
    value: IIF(count(healthCheck:responseid) > 0, IIF(average(SCORE(healthCheck:Q2)) >= 9, "Safe", IIF(average(SCORE(healthCheck:Q2)) >= 5, "Medium", "High")), "Unknown")
  }

  variable singleChoice #ooo {
    label: "oo"
    table: survey:
    option code {
      code: "Alert"
      score: 1
      label: "Alert"
    }
    option code {
      code: "Silent"
      score: 2
      label: "Silent"
    }
    value: IIF(survey:Q1 = "1", "Alert", IIF(IN(survey:status, "incomplete", "notanswered", "quotafull", "error", "screened"), "Silent"))

  }
}

config report #cr {
  paletteD: "#9BDC3E","#F6C54C","#EB666B","#E6E7E0"
  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Confirmit%20Demo/confirmit3Dlogo.jpg"
  palette: "#86ABE2","#4079D0","#1B6600","#2D9900","#9CCB00","#FEFE00","#F9BF00","#F18500","#EF6300","#F30000", "#AA0010", "#C0C0C0"
  paletteH: "#F6C54C","#E6E7E0","#9BDC3E","#EB666B"
  paletteM: "#E6E7E0","#9BDC3E","#F6C54C","#EB666B"
  formatter date #date11 {
    formatString: "DD MMM YYYY"
    emptyValue: "None"
  }
  formatter date #date12 {
    locale: en
    formatString: "DD MMM YYYY"
  }
  formatter date #month {
    locale: en
    formatString: "MMM YYYY"

  }
  formatter date #dateFormat {
    inputFormat: "YYYYMM"
    formatString: "MMMM"
  }

  formatter value #valueFMT {
    emptyValue: " "
  }
  formatter number #formatterID {
    numberDecimals: 0
    prefix: "$ "
    decimalSeparator: "."
    integerSeparator: " "
    shortForm: true
  }

  formatter number #formatterLTR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    emptyValue: "-"
  }
  formatter number #formatterRR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    postfix: " %"
  }

  formatter color #formatterColor {
    thresholds: #009900 >=9 , #b34700 >=7, #b30000 >=0
  }
  formatter color #formatterColor2 {
    thresholds: #0099AA >=9 , #b347AA >=7, #b300AA >=0
  }
  formatter number #metricFormat {
    numberDecimals: 1
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
  }

  formatter number #responsesFormat {
    numberDecimals: 0
    shortForm: false
  }

  formatter color #riskStringFormatter {
    thresholds: Unknown = 0 , Low = 1, Medium = 2, High = 3
  }

  formatter color #valueCases {
    thresholds: #ff0000 >=1, #31363e >=0
  }
  formatter color #backgroundColorFormatter {
    thresholds: #e8f8e0 >= 8.5, #ffeed6 >= 6.5, #fedfe2 >= 0
  }
  formatter color #valueColorFormatter {
    thresholds: #5ba35d >= 8.5, #ffa156 >= 6.5, #dd3435 >= 0
  }

  formatter date #dateForm {
    inputFormat: "YYYYMM"
    formatString: "MMM YY"
  }
}
layoutArea toolbar {
  filter multiselect {
    label: "DV"
    option checkbox {
      value: accounts:oo = "Safe"
      label: "Safe"
    }
    option checkbox {
      value: accounts:oo = "Medium"
      label: "Medium"
    }
    option checkbox {
      value: accounts:oo = "High"
      label: "High risk"
    }
  }
  filter multiselect #accountOwenr {
    label: "Account Owner"
    optionsFrom: accounts:AccountOwner
  }
  filter multiselect #risk {
    label: "Revenue Risk"
    filterType: postAggregate
    option checkbox #a {
      label: "High"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10
    }
    option checkbox #b {
      label: "Medium"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(surveyR:respid) * 100 > 4 AND average(SCORE(survey:Q1)) < 7 OR average(SCORE(healthCheck:NPS)) < 5
    }
    option checkbox #c {
      label: "Low"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(surveyR:respid) * 100 > 4 AND average(SCORE(survey:Q1)) > 6 AND count(healthCheck:responseid) > 0 AND average(SCORE(healthCheck:NPS)) > 6 OR count(healthCheck:responseid) > 0
    }

  }

  filter multiselect #region {
    label: "Region"
    optionsFrom: accounts:SalesRegion
  }

  filter multiselect #role {
    label: "Role"
    option checkbox #r1 {
      label: "Decision maker"
      value: contacts:contactRole = "Decision maker"
    }
    option checkbox #r2 {
      label: "Influencer"
      value: contacts:contactRole = "Influencer"
    }

  }
  filter multiselect #period {
    label: "Reporting period"
    option checkbox #s1 {
      label: "Last quarter"
      value: survey:interview_start > 2017-09-30 AND survey:interview_start < 2018-01-01
    }
    option checkbox #s2 {
      label: "Last 6 months"
      value: survey:interview_start > 2017-10-23
    }
    option checkbox #s3 {
      label: "Last 12 months"
      value: survey:interview_start > 2017-01-23
    }

  }


  filter multiselect #renewal {
    label: "Renewal period"
    option checkbox #q1 {
      label: "Q1 2018"
      value: accounts:RenewalDate > 2018-01-01 AND accounts:RenewalDate < 2018-04-01
    }
    option checkbox #q2 {
      label: "Q2 2018"
      value: accounts:RenewalDate > 2018-03-31 AND accounts:RenewalDate < 2018-07-01
    }
    option checkbox #q3 {
      label: "Q3 2018"
      value: accounts:RenewalDate > 2018-06-30 AND accounts:RenewalDate < 2018-10-01
    }
    option checkbox #q4 {
      label: "Q4 2018"
      value: accounts:RenewalDate > 2018-09-30 AND accounts:RenewalDate < 2019-01-01
    }
  }
}

page #Accounts {
  label: "Accounts"

  widget portfolioBreakdown #REX {
    label: "Risk with DV"
    size: medium
    category: IIF(accounts:RenewalDate >= 2018-06-01, CalendarMONTH(accounts:RenewalDate))
    categoryFormat: dateForm
    segment: accounts:oo
    value: count(survey:responseid)
    palette: @cr.paletteD
  }

  widget portfolioBreakdown #R {
    label: "Portfolio Risk Assessment"
    size: small
    category: CalendarMONTH(accounts:RenewalDate)
    categoryFormat: dateForm
    segment: IIF(count(healthCheck:responseid, true, accounts:) > 0, IIF(average(SCORE(healthCheck:Q2), true, accounts:) >= 9, "Safe", IIF(average(SCORE(healthCheck:Q2), true, accounts:) >= 5, "Medium", "High")), "Unknown")
    value: count(survey:responseid)
    palette: @cr.paletteM
  }
  widget accountList {
    label: "Accounts"
    table: accounts:
    sortColumn: accountName1
    sortOrder: descending

    column value #accountName1 {
      label: "Name"
      value: accounts:AccountName
    }
  }
  widget recentResponses #yy {
    label: "yy"

    showHeader: true
    view comment #fff {
      lines: 4
    }
    view metric #metrics {
      valueColorFormatter: valueColorFormatter
      fontSize: large
      backgroundColorFormatter: transparent
    }
    size: medium
    table: survey:
    column response #x1 {
      sortBy: footer
      footer: survey:interview_end
      header: survey:FirstName + " " + survey:LastName + " - " + accounts:AccountName
      comment: survey:Q2
    }
    column metric #ltr2 {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      target: 10
      view: metrics
    }
  }
  widget topAccounts {
    table: accounts:
    size: small
    sortColumn: main
    navigateTo: Accountdetails
    hierarchy: accounts:ParentAccountID


    view metricWithChange #metrics {
      valueColorFormatter: valueColorFormatter
      fontSize: medium
    }

    column accounts #main {
      accountName: accounts:AccountName
      revenue: accounts:AnnualAccountValue

      value: accounts:AnnualAccountValue
    }

    column metric #ltr {
      value: average(score(survey:Q1))
      previous: average(score(survey:Q3))
      format: formatterLTR
      target: 10
      view: metrics
    }

  }
  widget kpi {
    label: "DV"
    tile kpi {
      value: SUM(accounts:NN)

    }
  }

}

page #AccountList {
  label: "Account List"

  widget accountList {
    table: accounts:
    label: "Accounts"
    sortColumn: openCases
    sortOrder: descending
    size: large
    navigateTo: ContactList
    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }
    hierarchy: accounts:ParentAccountID

    column hierarchy #accountName {
      label: "Account Name "
      value: accounts:AccountName
      rowHeader: true
    }

    column value {
      label: "Derived variable"
      value: accounts:oo
    }
    column value #accountMan {
      label: "Account Owner"
      value: accounts:AccountOwner
    }
    column value #risk {
      label: "Risk Level"
      value: IIF(average(SCORE(survey:Q1)) < 7, "H", IIF(average(SCORE(survey:Q1)) > 8, "L", IIF(COUNT(survey:responseid) < 1, "U", "M")))

    }
    column value #ltr {
      label: " LTR "
      value: average(SCORE(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }
    column value #oast {
      label: "OSAT"
      value: average(SCORE(survey:Q4))
      format: metricFormat
      view: metrics
    }
    column value #openCases {
      label: "Cases"
      value: COUNT(cases:CaseId)
    }
    column value #responses {
      label: "Responses"
      value: COUNT(survey:responseid, survey:status = "complete")
      sortable: true
      align: center
    }
    column value #rate {
      label: "Response Rate"
      value: COUNT(survey:responseid, survey:status = "Complete") * 100 / COUNT(survey:respid)
      format: formatterRR
      sortable: true
      align: center
    }
    column value #noResp {
      label: "No Response"
      value: COUNT(survey:responseid) - COUNT(survey:responseid, survey:status = "Complete")
      sortable: true
      align: center
    }

  }
}

page #ContactList {
  label: "Contact List"

  widget contactList #hg {
    table: survey:
    label: "Contacts"
    inHierarchy: accounts:ParentAccountID
    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    column value #accountNN {
      label: "Company"
      value: survey:AccountName
    }

    column value #firstName {
      label: "First Name"
      value: survey:FirstName
    }

    column value #lastName {
      label: "Last Name"
      value: survey:LastName
    }
    column value #role {
      label: "Role"
      value: survey:ContactRole
    }

    column value #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: metricFormat
      view: metrics
    }
    column value #openCases {
      label: "Cases"
      value: COUNT(cases:CaseId)
    }

    column value #lastResponse {
      label: "Last response"
      value: max(survey:interview_end)
      format: date11
    }


    column value #comments {
      label: "Comments"
      value: MAX(survey:Q2, survey:interview_start = max(survey:interview_start))
    }
    column value #commentsN {
      label: "Value of comments"
      value: COUNT(survey:Q2)
    }

  }

}


page #Start {
  label: "Start"

  widget portfolioBreakdown {
    label: "Business vs Satisfaction"
    size: large
    category: survey:Industry
    segment: survey:Q1
    value: count(survey:responseId)
    percent: on
    //palette: @cr.palette
    format: formatterLTR
    navigateTo: AccountList
  }
}

page #Datebreakdown {
  label: "Date breakdown"

  widget portfolioBreakdown {

    label: "Month vs Satisfaction"
    size: large

    category: CalendarMonth(accounts:RenewalDate)
    segment: IIF(count(healthCheck:responseid, true, accounts:) > 0, IIF(average(SCORE(healthCheck:Q2), true, accounts:) >= 9, 1, IIF(average(SCORE(healthCheck:Q2), true, accounts:) >= 5, 2, 3)), 0)

    value: count(survey:responseId)
    format: floatNumber

    categoryFormat: dateFormat
    palette: @cr.palette
    navigateTo: LoneCuts
  }

  widget portfolioBreakdown #portfolioBreakdownWidget_2 {

    label: "Month vs Satisfaction (percent)"
    size: large

    category: Year(survey:interview_start)
    segment: survey:Q1
    value: count(survey:responseId)
    percent: on

    palette: @cr.palette
  }
}

page #LoneCuts {
  label: "Lone Cuts"

  widget portfolioBreakdown {
    label: "Q1 trend"
    size: large

    category: calendarMonth(survey:interview_start)
    categoryFormat: dateFormat
    value: average(score(survey:Q1))
    format: formatterLTR

  }

  widget portfolioBreakdown #portfolioBreakdownWidget_2 {
    label: "Responses per year (segments)"
    size: large

    segment: year(survey:interview_start)

    value: count(survey:responseid)
    percent: on
    navigateTo: AccountList
  }
  widget portfolioBreakdown #z1 {
    label: "Case Management Risk"
    size: small
    category: Year(survey:interview_start)
    segment: survey:ooo
    value: count(survey:)
  }
}

title "Artu Demo report"
//Do not edit please

config hub {

  hub: 101354
  table accounts = crmdata.ArtuAccountHierarchy //crmdata.externalAccounts   //p1028432.respondent
  table accounts2 = crmdata.externalAccounts // workaround for fetching data that are set to be Categorical
  table survey = p1863845164.response  //p1027835.response
  table contacts = p1864143727.response //p1028592.response
  table healthCheck = p1863840407.response //p1028039.response
  table cases = am.CASE
  table respondent = p1863845164.respondent //p1027835.respondent
  table revenue = crmdata.Historical_Revenue


  relation oneToMany #rel1 {
    primaryKey: accounts:AccountID
    foreignKey: contacts:AccountID
  }
  relation oneToMany #rel2 {
    primaryKey: accounts:AccountID
    foreignKey: healthCheck:AccountID
  }
  relation oneToMany #rel3 {
    primaryKey: accounts:AccountID
    foreignKey: revenue:AccountID
  }
  relation oneToOne #rel4 {
    primaryKey: accounts2:AccountID
    foreignKey: accounts:AccountID
  }
}

custom properties #cp {
  npsTarget: 50
  osatTarget: 9
  completeSurv: COUNT(survey:responseid, survey:status = "Complete")
  ltrValue: average(score(survey:Q1))
  ltrTarget: 8
  healthTarget: 8
  revenueDiff: (accounts:AnnualAccountValue - sum(revenue:AnnualAccountValue, revenue:Year = 2015)) / accounts:AnnualAccountValue * 100
  revenueRiskValue: IIF(@cp.revenueDiff < -10, 3, IIF(@cp.revenueDiff < 10, 2, 1))
  renewalRiskValue: IIF(@cp.rateValue < 5, 0, IIF(@cp.ltrValue < 7 AND average(SCORE(healthCheck:Renew)) < 7, 3, IIF(@cp.ltrValue > 6 AND average(SCORE(healthCheck:Renew)) > 6, 1, 2)))
  renewalRiskText: IIF(@cp.renewalRiskValue = 0, "Unknown", IIF(@cp.renewalRiskValue = 3, "High", IIF(@cp.renewalRiskValue = 1, "Low", "Medium")))
  risk1: (average(SCORE(healthCheck:NPS)) + average(SCORE(healthCheck:Renew)) + average(SCORE(healthCheck:OSAT))) / 3
  risk3: IIF(average(SCORE(survey:Q1)) < 7, "H!", IIF(average(SCORE(survey:Q1)) > 8, "L", IIF(COUNT(survey:responseid) < 1, "U", "M")))
  risk4: IIF(COUNT(survey:responseid, survey:status = "complete") / COUNT(survey:responseid) < 0.05, "Unknown", IIF(average(SCORE(survey:Q1)) < 7 AND average(SCORE(healthCheck:Renew)) < 7, "High", IIF(average(SCORE(survey:Q1)) > 6 AND average(SCORE(healthCheck:Renew)) > 6, "Safe", "Medium")))
  riskLogo: IIF(average(SCORE(survey:Q1)) < 7, @cp.highRiskLogo, IIF(average(SCORE(survey:Q1)) > 8, @cp.blankLogo, IIF(COUNT(survey:responseid) < 1, @cp.blankLogo, @cp.warningLogo)))
  riskValue: @cp.revenueRiskValue
  riskTarget: 10
  rateInvites: COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
  rateResponses: @cp.completeSurv
  rateValue: @cp.rateResponses / @cp.rateInvites * 100
  casesValue: COUNT(cases:CaseId, cases:SystemStatus = "Open")
  fullContactName: contacts:FirstName + " " + contacts:LastName
  currentPeriod: healthCheck:interview_start > 2016-06-22
  previousPeriod: healthCheck:interview_start <= 2016-06-22
  highRiskLogo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/autumnblaze.png"
  warningLogo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/tangerinedream.png"
  blankLogo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/transparent.png"
  contactLogo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/mch/53633418-5037-4CEB-AF68-D8616D95094B.jpg"
  currentPeriodFilter: survey:interview_start > 2016-01-01
  previousPeriodFilter: survey:interview_start <= 2016-01-01
}

config report #cr {
  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/artu-logo.png"
  formatter number #formatterLTR {
    numberDecimals: 2
    decimalSeparator: "."
  }
  formatter number #formatterRR {
    numberDecimals: 0
    decimalSeparator: "."
    postfix: "%"
  }
  formatter number #customEmpty {
    numberDecimals: 0
    emptyValue: "-"
  }
  formatter number #currency {
    numberDecimals: 0
    prefix: "$ "
    decimalSeparator: "."
    integerSeparator: " "
    shortForm: true
  }
  formatter objectProperty #textPicker {
    property: text
  }
  formatter color #backgroundColor {
    thresholds: #e8f8e0 >= 8, #ffeed6 >= 6, #fedfe2 >= 0
  }
  formatter color #valueColor {
    thresholds: #388e3c >= 8, #ff6d00 >= 6, #d40000 >= 0
  }
  formatter date #DDMMMYYYY {
    format: "DD MMM YYYY"
    shortForm: true
    emptyValue: "-"
  }
  formatter date #dateRelative {
    locale: en
    shortForm: false
    relative: true
  }
  formatter text #commentFormat {
    useDots: true
    length: 68
    emptyValue: "-"
  }
  formatter color #riskTextColorFormatter {
    thresholds: #FA5263 >= 3, #000000 < 3//#FFBD5B = 2, #82D854 = 1 //, #E1EEE8 = 0
  }
  formatter color #riskTextBgColorFormatter {
    thresholds: rgba(0, 0, 0, 0) >= 0 //, #000000 < 3//#FFBD5B = 2, #82D854 = 1 //, #E1EEE8 = 0
  }
  formatter color #riskBgColorFormatter {
    thresholds: #FA5263 = 3, #FFBD5B = 2, #82D854 = 1 , #E1EEE8 = 0
  }
  formatter color #riskStringFormatter {
    thresholds: Unknown = 0 , Low = 1, Medium = 2, High = 3
  }
  formatter color #kpiColorFormatter {
    thresholds: #82D854 >= 100%, #FFBD5B >= 80%, #FA5263 < 80%
  }
}

layoutArea toolbar {
  filter multiselect {
    optionsFrom: survey:NPSSegment
  }
  filter multiselect {
    label: "Account Rating"
    option checkbox {
      label: "Gold"
      value: accounts:TotalAccountValue > 200000
    }
    option checkbox {
      label: "Silver"
      value: accounts:TotalAccountValue > 99999 AND accounts:TotalAccountValue < 199999
    }
    option checkbox {
      label: "Bronze"
      value: accounts:TotalAccountValue < 100000
    }
  }

  filter multiselect {
    optionsFrom: revenue:Year
  }
  filter singleselect #rp {
    label: "Reporting Period"
    global: false
    option radio {
      selected: true
      label: "Rolling Year"
      value: InYear(survey:interview_start, -1, 0, 2016-01-01)
      previous: InYear(survey:interview_start, -2, -1, 2016-01-01)
    }
    option radio {
      label: "Rolling Quarter"
      value: InQuarter(survey:interview_start, -1, 0, 2016-07-01)
      previous: InQuarter(survey:interview_start, -2, -1, 2016-07-01)
    }
    option radio {
      label: "Rolling Month"
      value: InMonth(survey:interview_start, -1, 0, 2016-07-01)
      previous: InMonth(survey:interview_start, -2, -1, 2016-07-01)
    }
  }
}



page #Overview {
  label: "Overview"


  widget kpi {
    label: "NPS"
    size: small
    tile kpi {
      label: "NPS"
      value: NPS(survey:Q1) * 100
      target: @cp.npsTarget
      min: -100
      max: 100
      format: formatterLTR
      targetFormat: formatterLTR
      gaugeColorFormat: kpiColorFormatter  // valueColor
      tile value {
        label: "Responses"
        value: count(survey:Q1, @cp.currentPeriodFilter)
        max: count(survey:responseid, @cp.currentPeriodFilter)
        format: integer
      }
      tile value {
        label: "Yearly change"
        value: average(score(survey:Q1), @cp.currentPeriodFilter) - average(score(survey:Q1), @cp.previousPeriodFilter)
        format: formatterLTR
      }
    }
  }
  widget kpi {
    label: "Overall Satisfaction"
    size: small
    tile kpi {
      label: "AVG"
      value: average(score(survey:Q4))
      target: @cp.osatTarget
      min: 0
      max: 10
      format: formatterLTR
      targetFormat: formatterLTR
      gaugeColorFormat: kpiColorFormatter       //valueColor
      tile value {
        label: "Responses"
        value: count(survey:responseid, survey:status = "Complete")// AND @cp.currentPeriodFilter)
        max: count(survey:responseid, @cp.currentPeriodFilter)
        format: integer
      }
      tile value {
        label: "Yearly change"
        value: average(score(survey:Q4), @cp.currentPeriodFilter) - average(score(survey:Q4), @cp.previousPeriodFilter)
        format: formatterLTR
      }
    }
  }
  widget portfolioBreakdown {
    label: "Portfolio Breakdown by Role"
    size: small

    category: contacts:ContactRole
    segment: survey:NPSSegment
    value: count(survey:responseId)

    percent: on
  }

  widget portfolioBreakdown #z {
    info: "asdfuasdlkjfhalsdjkfhalskdjfh"
     //May07 NSA: colous are messed up, wong colours sematics: safe is red, shoould be green
    label: "Accounts Risk Groups"
    size: small
    category: accounts:RenewalYear
    segment: IIF(count(healthCheck:responseid, true, accounts:) > 0, IIF(average(SCORE(healthCheck:Renew), true, accounts:) >= 9, "Safe", IIF(average(SCORE(healthCheck:Renew), true, accounts:) >= 5, "Medium", "High")), "Unknown")
    value: count(survey:responseid)  //((sum(revenue:AnnualRevenue, revenue:year=2017))
    navigateTo: Accounts
  }

  widget portfolioBreakdown #rev {
    label: "Revenue Risk Assessment"
    size: small
    category: CalendarMONTH(accounts:RenewalDate)
    segment: IIF(count(healthCheck:responseid, true, accounts:) > 0, IIF(average(SCORE(healthCheck:Renew), true, accounts:) >= 9, "Safe", IIF(average(SCORE(healthCheck:Renew), true, accounts:) >= 5, "Medium", "High")), "Unknown")
    value: sum(accounts:TotalAccountValue)
    format: currency
  }
  widget recentResponses #IV {
    label: "Account Manager View"
    table: healthCheck:
    size: small
    navigateTo: Account
    lines: 3
    view metric #metrics {
      valueColorFormatter: valueColor
      fontSize: large
      backgroundColorFormatter: transparent
    }
    column response {
      sortBy: footer
      footer: healthCheck:interview_end
      header: accounts:AccountName  //(AnswerText(accounts:AccountOwner) + " - ") + AnswerText(accounts:SalesRegion)
      comment: accounts:AccountOwner

    }
    column metric #ltr3 {
      label: "LTR estimate"
      value: average(score(healthCheck:NPS))
      target: 9
      view: metrics
    }
  }
  widget recentResponses #yy1 {
    label: "Customer Responses"
    showHeader: true
    navigateTo: Responseview
    view comment #fff {
      lines: 3
    }
    view metric #metrics {
      valueColorFormatter: valueColor
      fontSize: large
      backgroundColorFormatter: transparent
    }
    size: small
    table: survey:
    column response #x11 {
      sortBy: footer
      footer: survey:interview_end
      header: survey:FirstName + " " + survey:LastName + " - " + accounts:AccountName
      comment: survey:Q2
      commentFormat: commentFormat
    }
    column metric #ltr2 {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      target: 10
      view: metrics
    }
  }

  widget topAccounts {
    table: accounts:
    size: small
    sortColumn: main
    navigateTo: Account
    hierarchy: accounts:ParentAccountID
    view metricWithChange #metrics {
      valueColorFormatter: valueColor
      fontSize: medium
    }
    column accounts #main {
      accountName: accounts:AccountName
      revenue: accounts:AnnualAccountValue
      value: accounts:AnnualAccountValue
    }
    column metric #ltr {
      value: average(score(survey:Q1), @cp.currentPeriodFilter)
      previous: average(score(survey:Q1), @cp.previousPeriodFilter)
      format: formatterLTR
      target: @cp.ltrTarget
      view: metrics
    }
  }
}



page #Accounts {
  label: "Accounts"


  widget search {
    layoutArea: "header"    // not required ("header" by default)
    source search #source1_id {
      table: accounts //the name of the table in hub config (this is the table we search through)
      value: accounts:AccountName + " - " + accounts:AccountId //either field or fields-expression to search by
      navigateTo: Account //the name of the page to navigate when an item is clicked in the search suggestion
      iconType: "account"
    }
  }

  widget accountList {
    label: "Accounts"
    size: large
    table: accounts:
    sortColumn: accountName
    sortOrder: ascending
    navigateTo: Account
    hierarchy: accounts:ParentAccountID
  // views
    view metricWithChange #metrics {
      backgroundColorFormatter: backgroundColor
      valueColorFormatter: valueColor
      fontSize: small
    // roundCorners:true
    }
    view metric #risk {
      backgroundColorFormatter: riskTextBgColorFormatter
      valueColorFormatter: riskTextColorFormatter
      fontSize: small

    // roundCorners:true
    }

  // columns
    column hierarchy #accountName {
      label: "Accounts"
      value: accounts:AccountName
      rowHeader: true
    }

    column metric #revenueRisk {
      label: "Revenue Risk"
      value: @cp.riskValue
      target: 1
      format: riskStringFormatter
      valueColorFormatter: riskBgColorFormatter
      //view: iconSmall
      view: risk
    }
    column metric #renewalRisk {
      label: "Renewal Risk"
      value: @cp.renewalRiskValue
      target: 1
      format: riskStringFormatter
      //view: iconSmall
      view: risk
    }
    column metric #LTR {
      label: "LTR"
      value: average(score(survey:Q1), @rp.selectedOption.value)
      previous: average(score(survey:Q1), @rp.selectedOption.previous)
      target: @cp.ltrTarget
      format: formatterLTR
      align: left
      view: metrics
    }

    column metric #osat {
      label: "OSAT"
      value: average(score(survey:Q4), @cp.currentPeriodFilter)
      previous: average(score(survey:Q4), @cp.previousPeriodFilter)
      format: formatterLTR
      view: metrics
      target: @cp.osatTarget
      align: left
    }
    column metric #health11 {
      label: "Internal View"
      value: average(score(healthCheck:Renew), @cp.currentPeriod)
      previous: average(score(healthCheck:Renew), @cp.previousPeriod)
      target: @cp.healthTarget
      format: formatterLTR
      view: metrics
      align: left
    }
    column value #total {
      label: "Revenue ($)"
      value: accounts:TotalAccountValue
      format: currency
    }
    column value #case1 {
      label: "Cases"
      value: @cp.casesValue
      format: customEmpty
    }

    column value #responses {
      label: "Responses"
      value: @cp.completeSurv
      align: right
    }
    column value #rate {
      label: "Response Rate"
      value: @cp.rateValue
      format: formatterRR
    }
    column value #noResp {
      label: "No Response"
      align: right
      value: COUNT(survey:responseid) - @cp.completeSurv //COUNT(survey:responseid,survey:smtpstatus="Sent")
    }
    column value #survCount {
      label: "Surveys"
      value: count(survey:responseid)
      align: right
    }
  }
}

page account #Account {
  label: "Account"

  widget search {
    table: accounts:
    layoutArea: "header"
    value: accounts:AccountName + " - " + accounts:AccountId
    navigateTo: AccountPage
    iconType: "account"
  }
  widget title {
    table: accounts:
    layout column {
      tile value #c {
        value: accounts:AccountName
      }
    }
  }
  widget summary {
    table: accounts:
    hierarchy: accounts:ParentAccountID
    size: large
    tile metric {
      label: "LTR Avg"
      value: @cp.ltrValue
      target: @cp.ltrTarget
    }
    tile metric {
      label: "Account Manager View"
      value: average(score(healthCheck:Renew))
      target: @cp.healthTarget
    }
    tile risk {
      label: "Renewal Risk"
      value: @cp.renewalRiskValue
      target: 9
      min: 1
      max: 3
      renewal: accounts:renewalDate
      revenue: accounts:TotalAccountValue
      textValue: @cp.renewalRiskText
      format: valueFormatter
      backgroundColorFormatter: riskBgColorFormatter
    }
    tile responseRate {
      invites: @cp.rateInvites
      responses: @cp.rateResponses
    }
    tile casesStatus {
      open: @cp.casesValue
      overdue: 0
    }
  }

  widget contactList #hg {
    label: "Contacts"
    table: contacts:
    size: large
    sortColumn: name
    sortOrder: descending
    navigateTo: Contact
    view metricWithChange #metrics {
      backgroundColorFormatter: backgroundColor
      valueColorFormatter: valueColor
      fontSize: small
    }
    column value #name {
      label: "Name"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #company {
      label: "Company"
      value: contacts:AccountName
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }
    column metric #LTR {
      label: "LTR"
      value: average(score(survey:Q1), @cp.currentPeriodFilter)
      previous: average(score(survey:Q1), @cp.previousPeriodFilter)
      target: @cp.ltrTarget
      format: formatterLTR
      align: left
      view: metrics
    }

    column metric #osat {
      label: "OSAT"
      value: average(score(survey:Q4), @cp.currentPeriodFilter)
      previous: average(score(survey:Q4), @cp.previousPeriodFilter)
      format: formatterLTR
      view: metrics
      target: @cp.osatTarget
      align: left
    }
    column value #openCases {
      label: "Cases"
      value: @cp.casesValue
    }
    column value #lastResponse {
      label: "Last response"
      value: Year(max(survey:interview_end))
      asign: center
    }
    column value #comments {
      label: "Comments"
      value: LAST(survey:Q2, survey:interview_start, survey:interview_start > 2006-01-01)  //survey:NPSSegment='passive')  //, survey:interview_start, COUNT(cases:CaseId) > 0)
    }

  }
  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: datecreated
    sortOrder: descending

    view link #openLink {
      label: "View Case"
    }

    column value #datecreated {
      label: "Created"
      value: cases:DateCreated
      asign: center
      format: dateRelative
    }
    column value #dueDate {
      label: "Due"
      value: cases:DateDue
      asign: center
      format: dateRelative
    }
    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000920", "Technology issue", "NPS Detractors"))
    }
    column value #issueCat {
      label: "Issue Category"
      value: cases:lk_2906
      format: textPicker
    }
    column value #res {
      label: "Resolution"
      value: cases:lk_2907
      format: textPicker
    }
    column value #f {
      label: "CaseLink "
      value: cases:CaseLink
      view: openLink
    }
  }
}

page contact #Contact {
  label: "Contact"

  widget search {
    table: contacts:
    layoutArea: "header"
    value: @cp.fullContactName
    navigateTo: ContactList
  }
  widget title {
    table: contacts:
    layout column {
      tile icon {
        value: @cr.logo
      }
    }
    layout column {
      layout row {
        tile value {
          value: contacts:FirstName + " " + contacts:LastName
        }
        tile role {
          value: contacts:ContactRole
        }
      }
      layout row {
        tile company {
          value: contacts:AccountName
        }
      }
    }
  }

  widget summary {
    size: large
    table: contacts:
    tile contactDetails #cc {
      email: contacts:email
      title: contacts:AccountName
      phone: contacts:Phone
      role: contacts:ContactRole
      industry: contacts:Industry
    }
    tile accountDetails #cc4 {
      accountOwner: accounts2:AccountOwnerManager //+ " (") + (accounts:AccountOwnerManagerEmail + ")")
      salesManager: accounts2:SalesLeader1
      region: accounts2:WorldRegion
      revenue: accounts:AnnualAccountValue
      renewalDate: accounts:RenewalDate
    }
    tile metric {
      label: "LTR"
      value: @cp.ltrValue
      target: @cp.ltrTarget
    }

    tile surveyResponses #da {
      label: "Survey Responses"
      total: count(survey:responseid)
      completed: @cp.completeSurv
    }
  }

  widget contactSurveys {
    label: "Surveys"
    table: survey:
    sortColumn: is
    size: large
    sortOrder: descending
    navigateTo: Responseview

    view metricWithChange #metrics {
      backgroundColorFormatter: backgroundColor
      valueColorFormatter: valueColor
      fontSize: small
    }

    column value #s2 {
      label: "Status"
      value: survey:status
    }

    column value #is {
      label: "Date"
      value: survey:interview_start
      format: dateRelative
    }

    column metric #s3 {
      label: "LTR"
      value: average(score(survey:Q1), @cp.currentPeriodFilter)
      target: @cp.ltrTarget
      format: formatterLTR
      align: left
      view: metrics

    }
    column metric #osat {
      label: "OSAT"
      value: average(score(survey:Q4), @cp.currentPeriodFilter)
      format: formatterLTR
      view: metrics
      target: @cp.osatTarget
      align: left
    }

    column value #s6 {
      label: "Comments"
      value: survey:Q8
    }
  }
}

page account #Responseview {
  label: "Response view"

  widget contactSurveyResponse {
    view title #defaultSurveyResponseTitle {
    }


    size: medium
    surveyResponseTitle {

      tile title #rt {
        value: contacts:FirstName + " " + contacts:LastName + " - Relationship Survey"
        surveyName: survey:responseid
        view: defaultSurveyResponseTitle
      }
    }
    summary {
      rows: 4

      tile list #list1 {

        item value {
          value: survey:UploadedDate
          label: "Received"
          format: DDMMMYYYY
        }
        item value {
          value: survey:status
          label: "Status"
        }
        item email {
          value: survey:interview_start
          label: "Interview Start"
        }
        item value {
          value: survey:interview_end
          label: "Interview End"
        }
      }
      tile list #list2 {
        item value {
          value: "Relationship Survey"
          label: "Source"
        }
        item email {
          value: survey:responseid
          label: "Response ID"
        }
        item value {
          value: contacts:contactid
          label: "Respondent ID"
        }
      }
    }

    tab {
      label: "All"
      tile list {
        label: " "
        item comment {
          label: "First Name"
          value: contacts:FirstName
        }
        item comment {
          label: "Last Name"
          value: contacts:LastName
        }
        item comment {
          label: "Company name"
          value: accounts:AccountName
        }
        item comment {
          label: "Title"
          value: contacts:Title
        }
        item comment {
          label: "Role"
          value: contacts:ContactRole
        }
        view: defaulViewForListTile
      }
      tile list {
        label: "Key Metrics"
        item bar {
          label: "Likelihood to Recommend"
          value: average(score(survey:Q1))
        }
        item bar {
          label: "Overall Satisfaction"
          value: average(score(survey:Q4))
        }
        item comment {
          label: "Satisfaction with Technology"
          value: survey:Q8
        }
        view: defaulViewForListTile
      }
      tile list {
        label: "Product Satisfaction"
        item bar {
          label: "Technology"
          value: average(score(survey:Q7))
        }
        item bar {
          label: "Product is scalable"
          value: average(score(survey:Q9.1))
        }
        item bar {
          label: "Product is easy to use"
          value: average(score(survey:Q9.2))
        }
        item bar {
          label: "Product delivers results"
          value: average(score(survey:Q9.3))
        }
        view: defaulViewForListTile
      }
      tile list {
        label: "Service Satisfaction"
        item bar {
          label: "Provide Added Value"
          value: average(score(survey:Q3))
        }
        item bar {
          label: "Support business needs"
          value: average(score(survey:Q12))
        }
        view: defaulViewForListTile
      }
    }
    tab {
      label: "Comments"
      tile list {
        label: "Key"
        item comment {
          label: "label1"
          value: survey:Q2
        }
        item comment {
          label: "label2"
          value: survey:Q6
        }
      }
      view: defaulViewForListTile
    }
    tab {
      label: "CASE DATA"
      tile list {
        label: "NPS Detractor Alert"
        item bar {
          label: "Likelihood to Recommend"
          value: average(score(survey:Q1))
        }
        item bar {
          label: "Overall Satisfaction"
          value: average(score(survey:Q4))
        }
        item comment {
          label: "Satisfaction with Technology"
          value: survey:Q8
        }
        view: defaulViewForListTile
      }
      tile list {
        label: "Product Satisfaction"
        item bar {
          label: "Technology"
          value: average(score(survey:Q7))
        }
        item bar {
          label: "Product is scalable"
          value: average(score(survey:Q9.1))
        }
        item bar {
          label: "Product is easy to use"
          value: average(score(survey:Q9.2))
        }
        item bar {
          label: "Product delivers results"
          value: average(score(survey:Q9.3))
        }
        view: defaulViewForListTile
      }
      tile list {
        label: "Service Satisfaction"
        item bar {
          label: "Provide Added Value"
          value: average(score(survey:Q3))
        }
        item bar {
          label: "Support business needs"
          value: average(score(survey:Q12))
        }
        view: defaulViewForListTile
      }
    }
  }
}
title "Terry's risk report"

//NSA 20Jan : updated risk model (not final) and cosmetic changes applied to case table and Contact Title added some come
config access {
  portalid: 1870
  ssoConfig: Confirmit_Salesforce
}

config hub {
  hub: 14900
  table accounts = custom.Account_2      //accounts custom table
  table survey = p1850259384.response  //relationship survey
  table contacts = p1862934241.response
  table healthCheck = p1860215844.response      //healthcheck survey
  table cases = am.CASE
  table respondent = p1850259384.respondent
  table revenue = custom.Historical_Revenue  // historical revenue custom table.
  table new = custom.Account_2
  table ejournal = custom.eJournal

  //accounts --> revenue
  relation oneToMany #rel3 {
    primaryKey: accounts:accountID
    foreignKey: revenue:accountID
  }

  // accounts --> Health
  relation oneToMany #rel2 {
    primaryKey: accounts:AccountID
    foreignKey: healthCheck:shortAccountID

  }
  // accounts --> contact db --> survey
  relation oneToMany #rel4 {
    primaryKey: accounts:AccountID
    foreignKey: contacts:shortAccountID
  }
  //accounts --> eJournal
  relation oneToMany #rel5 {
    primaryKey: accounts:eJournalAccountNumber
    foreignKey: ejournal:compid
  }

}
layoutArea toolbar {

  filter multiselect #accountOwenr {
    label: "Account Owner"
    optionsFrom: accounts:AccountOwner
  }
  filter multiselect #risk {
    label: "Revenue Risk"
    filterType: postAggregate
    option checkbox #a {
      label: "High"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10
    }
    option checkbox #b {
      label: "Medium"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(respondent:respid) * 100 > 4 AND average(SCORE(survey:Q1)) < 7 OR average(SCORE(healthCheck:NPS)) < 5
    }
    option checkbox #c {
      label: "Low"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(respondent:respid) * 100 > 4 AND average(SCORE(survey:Q1)) > 6 AND count(healthCheck:responseid) > 0 AND average(SCORE(healthCheck:NPS)) > 6 OR count(healthCheck:responseid) > 0
    }

  }

  filter multiselect #region {
    label: "Region"
    optionsFrom: accounts:SalesRegion
  }

  filter multiselect #role {
    label: "Role"
    option checkbox #r1 {
      label: "Decision maker"
      value: contacts:contactRole = "Decision maker"
    }
    option checkbox #r2 {
      label: "Influencer"
      value: contacts:contactRole = "Influencer"
    }
  }
  filter multiselect #period {
    label: "Reporting period"
    option checkbox #s1 {
      label: "Last quarter"
      value: survey:interview_start > 2017-09-30 AND survey:interview_start < 2018-01-01
    }
    option checkbox #s2 {
      label: "Last 6 months"
      value: survey:interview_start > 2017-10-23
    }
    option checkbox #s3 {
      label: "Last 12 months"
      value: survey:interview_start > 2017-01-23
    }
  }

  filter multiselect #renewal {
    label: "Renewal period"
    option checkbox #q1 {
      label: "Q1 2018"
      value: accounts:RenewalDate > 2018-01-01 AND accounts:RenewalDate < 2018-04-01
    }
    option checkbox #q2 {
      label: "Q2 2018"
      value: accounts:RenewalDate > 2018-03-31 AND accounts:RenewalDate < 2018-07-01
    }
    option checkbox #q3 {
      label: "Q3 2018"
      value: accounts:RenewalDate > 2018-06-30 AND accounts:RenewalDate < 2018-10-01
    }
    option checkbox #q4 {
      label: "Q4 2018"
      value: accounts:RenewalDate > 2018-09-30 AND accounts:RenewalDate < 2019-01-01
    }
  }
}
custom properties #cp {
  // variables to be used by writing e.g. @cp.revenueRiskValue // cr =
  revenueRiskValue: IIF((sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10, 3, IIF((sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < 10, 2, 1))
}

config report #cr {
  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Confirmit%20Demo/confirmit3Dlogo.jpg"

  formatter date #date11 {
    shortForm: true
    emptyValue: "None"
  }
  formatter date #date12 {
    locale: en
    shortForm: false
  }
  formatter value #valueFMT {
    emptyValue: " "
  }
  formatter number #formatterID {
    numberDecimals: 0
    prefix: "$ "
    decimalSeparator: "."
    integerSeparator: " "
    shortForm: true
  }
  formatter number #formatterLTR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    emptyValue: "-"
  }
  formatter number #formatterRR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    postfix: " %"
  }

  formatter color #formatterColor {
    thresholds: #009900 >=9 , #b34700 >=7, #b30000 >=0
  }
  formatter color #formatterColor2 {
    thresholds: #0099AA >=9 , #b347AA >=7, #b300AA >=0
  }
  formatter number #metricFormat {
    numberDecimals: 1
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
  }

  formatter number #responsesFormat {
    numberDecimals: 0
    shortForm: false
  }

  formatter color #riskStringFormatter {
    thresholds: Unknown = 0 , Low = 1, Medium = 2, High = 3
  }

  formatter color #valueCases {
    thresholds: #ff0000 >=1, #31363e >=0
  }
  formatter color #backgroundColorFormatter {
    thresholds: #e8f8e0 >= 8.5, #ffeed6 >= 6.5, #fedfe2 >= 0
  }
  formatter color #valueColorFormatter {
    thresholds: #5ba35d >= 8.5, #ffa156 >= 6.5, #dd3435 >= 0
  }
  formatter objectProperty #textPicker {
    property: text
  }

  formatter color #riskColorFormatter {
    thresholds: #FA5263 >= 99%, #FFBD5B >=49%, #82D854 >0%
  }


}

page #AccountList {
  label: "Account List"

  widget markdown {
    size: medium

    markdown: "
## Confirmit Confidential Information"
  }
  widget accountList {
    label: "Accounts"
    table: accounts:
    sortColumn: healthrisk
    sortOrder: descending
    navigateTo: Account
    size: large

    hierarchy: accounts:ParentAccountID

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    column hierarchy #accountName {
      label: "Account Name "
      value: accounts:AccountName
      rowHeader: true
    }
    column value #accountMan {
      label: "Account Owner"
      value: accounts:AccountOwner
    }

    column value #healthrisk {
      label: "Health Risk"
      value: IIF(IIF(count(healthCheck:responseid) > 0, 1, 0) = 1, IIF(average(SCORE(healthCheck:Q2)) >= 9, 1, IIF(average(SCORE(healthCheck:Q2)) >= 5, 2, 3)), 0)
      align: center
      format: riskStringFormatter
    }

    column value #relrisk {
      label: "LTR Risk"
      value: IIF(COUNT(respondent:respid) = 0, 0, IIF(IIF(COUNT(survey:responseid, survey:status = "complete" OR survey:status = "incomplete") / COUNT(respondent:respid) * 100 < 5, 0, 1) = 1, IIF(average(SCORE(survey:Q1)) >= 9, 1, IIF(average(SCORE(survey:Q1)) > 6, 2, IIF(average(SCORE(survey:Q1)) > 0, 3, 0))), 0))
      align: center
      format: riskStringFormatter
    }

    column value #revRisk {
      label: "Revenue Risk "
      value: @cp.revenueRiskValue
      align: center
      format: riskStringFormatter
    }

    column metric #hh {
      label: "Health"
      value: average(score(healthCheck:Q2))
      format: formatterLTR
      view: metrics
      target: 9
    }
    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column value #rev2017 {
      label: "2017 rev"
      value: sum(revenue:AnnualRevenue, revenue:year = 2017)
      format: formatterID
      align: right
    }
    column value #rev2016 {
      label: "2016 rev"
      value: sum(revenue:AnnualRevenue, revenue:year = 2016)
      format: formatterID
      align: right
    }
    column value #revDiff {
      label: "Rev diff"
      value: sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)
      format: formatterID
      align: right
    }
    column value #revDiffPercentage {
      label: "Rev diff"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100
      format: formatterRR
      align: right
    }
    column value #tickets {
      label: "eJournal total"
      value: sum(ejournal:closedTickets)
    }
    column value #ticketsOpen {
      label: "eJournal Open"
      value: sum(ejournal:openTickets)
    }

    column value #case2 {
      label: "Cases"
      value: COUNT(cases:CaseId)
      align: center
      format: responsesFormat

    }
    column value #responses {
      label: "Responses "
      format: valueFMTnses
      value: COUNT(survey:responseid, survey:status = "complete" OR survey:status = "incomplete")
      align: center
    }
    column value #rate {
      label: "Response Rate"
      value: COUNT(survey:responseId, survey:status = "complete" OR survey:status = "incomplete") * 100 / COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
      format: formatterRR
      align: center
    }
    column value #noResp {
      label: "No Response"
      value: COUNT(respondent:respid, respondent:smtpstatus = "messagesent") - COUNT(survey:responseid, survey:status = "Complete")
      align: center
    }
  }
}

page account #Account {
  label: "Account"


  widget search {
    table: accounts:
    layoutArea: "header"
    value: accounts:AccountName + " " + accounts:AccountId
    navigateTo: AccountPage
    iconType: "account"
  }


  widget title {
    table: accounts:
    layout column {
      tile value #c {
        value: accounts:accountName
      }
    }
  }

  widget summary {
    size: large
    table: accounts:

    tile metric {
      label: "LTR Average"
      value: average(score(survey:Q1))
      target: 7
    }

    tile metric {
      label: "Account Owner View"
      value: average(score(healthCheck:Q1))
      target: 5
    }


    tile risk {
      label: "Revenue Risk"
        // need to tune formatting! add calculation
      value: @cp.revenueRiskValue
      textValue: IIF(@cp.revenueRiskValue = 3, "High", IIF(@cp.revenueRiskValue = 2, "Medium", IIF(@cp.revenueRiskValue = 1, "Low", "Unknown")))
      min: 1
      max: 3
      target: 0
      renewal: accounts:RenewalDate
      revenue: sum(revenue:AnnualRevenue, revenue:year = 2017)
      backgroundColorFormatter: riskColorFormatter
    }

    tile responseRate {
      invites: COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
      responses: COUNT(survey:responseId, survey:status = "complete" OR survey:status = "incomplete")
    }

    tile casesStatus {
      label: "Cases"
      open: COUNT(cases:CaseId)
      overdue: 0
    }
  }

  widget contactSurveys {
    label: "Internal View Survey"
    table: healthCheck:
    sortColumn: surveyDate
    sortOrder: ascending
    size: large

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    column value #accountMan {
      label: "Account Owner"
      value: accounts:AccountOwner
    }

    column date #surveyDate {
      label: "Date"
      value: healthCheck:interview_start
    }

    column metric #ltr {
      label: "LTR estimate"
      value: average(score(healthCheck:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column metric #ltr2 {
      label: "Renewal"
      value: average(score(healthCheck:Q2))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }
    column metric #ltr3 {
      label: "Growth Potential"
      value: average(score(healthCheck:Q5))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column metric #ltr4 {
      label: "Dependency on Services"
      value: average(score(healthCheck:Q11))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }
    column value #comments {
      label: "Comments: how to keep the customer"
      value: healthCheck:Q4
    }
  }

  widget contactList #hg {
    size: large
    label: "Account Contacts "
    table: contacts:
    sortColumn: name
    sortOrder: descending
    navigateTo: Contact
    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    view metric #ccc {
      valueColorFormatter: valueCases
    }
    column value #name {
      label: "Name"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #company {
      label: "Company"
      value: contacts:AccountName
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }

    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
    }
    column value #openCases {
      label: "Cases"
      value: COUNT(cases:CaseId)
      view: ccc
    }
    column value #lastResponse {
      label: "Last response "
      value: LAST(survey:interview_start, survey:interview_start)
      format: date11
      asign: center
    }
    column value #comments {
      label: "Comments"
      value: LAST(survey:Q2, survey:interview_start)
    }
  }

  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Date"
      value: cases:DateCreated
      align: center
      format: date12
    }

    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000818", "Health Check : At Risk", IIF(cases:Workflow = "1000819", "Health Check : High Potential", "Relationship : Recommend and/or Tech Detractors")))
    }
    column value #res {
      label: "Resolution"
      value: IIF(cases:lk_1548 = "5218" OR cases:lk_1548 = "5219" OR cases:lk_1548 = "5220", "Client specific", IIF(cases:lk_1548 = "5221" OR cases:lk_1548 = "5222" OR cases:lk_1548 = "5223", "Generic", IIF(cases:lk_1548 = "8319" OR cases:lk_1548 = "8320" OR cases:lk_1548 = "8321" OR cases:lk_1548 = "8322", "At risk: Action Taken", IIF(cases:lk_1548 = "8323" OR cases:lk_1548 = "8324", "High potential", "To Be Coded"))))
    }
    column value #link {

      label: "Action"
      value: cases:CaseLink
      view: link1
    }

  }
}

page contact #Contact {
  label: "Contact"


  widget search {
    table: contacts:
    layoutArea: "header"
    value: contacts:client_first_name + " " + contacts:client_last_name
    navigateTo: ContactList
  }

  widget title {
    table: contacts:
    layout column {
      tile icon {
        value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/magdalenas/defaultLogo.PNG"//"http://is1.mzstatic.com/image/thumb/Purple71/v4/89/51/f4/8951f4f1-fd6b-fa59-38b2-191140473b9a/source/175x175bb.jpg"
      }
    }
    layout column {
      layout row {
        tile value {
          value: contacts:FirstName + " " + contacts:LastName
        }
        tile role {
          value: contacts:ContactRole
        }
      }
      layout row {
        tile company {
          value: contacts:AccountName
        }
      }
    }
  }

  widget summary {
    size: large
    table: contacts:
    tile contactDetails #cc {
      title: contacts:Title
      role: contacts:ContactRole
      email: contacts:email
      phone: contacts:Phone
      industry: contacts:Industry
    }

    tile accountDetails #cc4 {
      accountOwner: contacts:AccountOwner
      salesManager: contacts:SalesLeader1
      region: contacts:WorldRegion
      revenue: contacts:AnnualAccountValue
      renewalDate: accounts:RenewalDate
      //rene
    }

    tile metric #a {
      label: "LTR"
      value: average(score(survey:Q1))
      target: 9
    }
    tile surveyResponses {
      total: count(respondent:respid)
      completed: count(survey:responseid, survey:status = "Complete")
    }
    tile casesStatus {
      label: Cases
      open: count(cases:CaseId)
      overdue: 0
    }
  }

  widget contactSurveys {
    label: "Surveys"
    table: survey:
    sortColumn: surveyDate
    sortOrder: ascending
    size: large

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
      //roundCorners:true
    }

    column value #status {
      label: "Status"
      value: survey:status
    }

    column date #surveyDate {
      label: "Date"
      value: survey:interview_end
    }

    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column value #case2 {
      label: "Cases"
      value: COUNT(cases:CaseId)
      align: center
      format: responsesFormat
    }

    column value #comments {
      label: "Comments"
      value: survey:Q2
    }
  }

  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending
    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Date"
      value: cases:DateCreated
      align: center
      format: date12
    }
    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000818", "Health Check : At Risk", IIF(cases:Workflow = "1000819", "Health Check : High Potential", "Relationship : Recommend and/or Tech Detractors")))
    }
    column value #res {
      label: "Resolution"
      value: IIF(cases:lk_1548 = "5218" OR cases:lk_1548 = "5219" OR cases:lk_1548 = "5220", "Client specific", IIF(cases:lk_1548 = "5221" OR cases:lk_1548 = "5222" OR cases:lk_1548 = "5223", "Generic", IIF(cases:lk_1548 = "8319" OR cases:lk_1548 = "8320" OR cases:lk_1548 = "8321" OR cases:lk_1548 = "8322", "At risk: Action Taken", IIF(cases:lk_1548 = "8323" OR cases:lk_1548 = "8324", "High potential", "To Be Coded"))))
    }
    column link #caseLink {
      label: "Case Link"
      value: cases:CaseLink
      view: link1
    }

  }
}
title "Terry's risk report"

//NSA 20Jan : updated risk model (not final) and cosmetic changes applied to case table and Contact Title added some come

config access {
  portalid: 1870
  ssoConfig: Confirmit_Salesforce
}

// workaround to avoid Compiler Error for config access block
config pulse

config hub {
  hub: 14900
  table accounts = custom.Account_2      //accounts custom table
  table survey = p1850259384.responseid  //relationship survey
  table contacts = p1862934241.responseid
  table healthCheck = p1860215844.responseid      //healthcheck survey
  table cases = am.CASE
  table respondent = p1850259384.respondent
  table revenue = custom.Historical_Revenue  // historical revenue custom table.
  table new = custom.Account_2
  table ejournal = custom.eJournal

  //accounts --> revenue
  relation oneToMany #rel3 {
    primaryKey: accounts:accountID
    foreignKey: revenue:accountID
  }

  // accounts --> Health
  relation oneToMany #rel2 {
    primaryKey: accounts:AccountID
    foreignKey: healthCheck:shortAccountID

  }
  // accounts --> contact db --> survey
  relation oneToMany #rel4 {
    primaryKey: accounts:AccountID
    foreignKey: contacts:shortAccountID
  }
  //accounts --> eJournal
  relation oneToMany #rel5 {
    primaryKey: accounts:eJournalAccountNumber
    foreignKey: ejournal:compid
  }

}
layoutArea toolbar {
  filter multiselect #accountOwenr {
    label: "Account Owner"
    optionsFrom: accounts:AccountOwner
  }
  filter multiselect #risk {
    label: "Revenue Risk"
    filterType: postAggregate
    option checkbox #a {
      label: "High"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10
    }
    option checkbox #b {
      label: "Medium"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(respondent:respid) * 100 > 4 AND average(SCORE(survey:Q1)) < 7 OR average(SCORE(healthCheck:NPS)) < 5
    }
    option checkbox #c {
      label: "Low"
      value: COUNT(survey:responseid, survey:status = "complete") / COUNT(respondent:respid) * 100 > 4 AND average(SCORE(survey:Q1)) > 6 AND count(healthCheck:responseid) > 0 AND average(SCORE(healthCheck:NPS)) > 6 OR count(healthCheck:responseid) > 0
    }

  }

  filter multiselect #region {
    label: "Region"
    optionsFrom: accounts:SalesRegion
  }

  filter multiselect #role {
    label: "Role"
    option checkbox #r1 {
      label: "Decision maker"
      value: contacts:contactRole = "Decision maker"
    }
    option checkbox #r2 {
      label: "Influencer"
      value: contacts:contactRole = "Influencer"
    }

  }
  filter multiselect #period {
    label: "Reporting period"
    option checkbox #s1 {
      label: "Last quarter"
      value: survey:interview_start > 2017-09-30 AND survey:interview_start < 2018-01-01
    }
    option checkbox #s2 {
      label: "Last 6 months"
      value: survey:interview_start > 2017-10-23
    }
    option checkbox #s3 {
      label: "Last 12 months"
      value: survey:interview_start > 2017-01-23
    }

  }


  filter multiselect #renewal {
    label: "Renewal period"
    option checkbox #q1 {
      label: "Q1 2018"
      value: accounts:RenewalDate > 2018-01-01 AND accounts:RenewalDate < 2018-04-01
    }
    option checkbox #q2 {
      label: "Q2 2018"
      value: accounts:RenewalDate > 2018-03-31 AND accounts:RenewalDate < 2018-07-01
    }
    option checkbox #q3 {
      label: "Q3 2018"
      value: accounts:RenewalDate > 2018-06-30 AND accounts:RenewalDate < 2018-10-01
    }
    option checkbox #q4 {
      label: "Q4 2018"
      value: accounts:RenewalDate > 2018-09-30 AND accounts:RenewalDate < 2019-01-01
    }
  }
}

custom properties #cp {
  // variables
  revenueRiskValue: IIF((sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < -10, 3, IIF((sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100 < 10, 2, 1))
}

config report {
  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Confirmit%20Demo/confirmit3Dlogo.jpg"

  formatter date #date11 {
    shortForm: true
    emptyValue: "None"
  }
  formatter date #date12 {
    locale: en
    shortForm: false
  }
  formatter value #valueFMT {
    emptyValue: " "
  }
  formatter number #formatterID {
    numberDecimals: 0
    prefix: "$ "
    decimalSeparator: "."
    integerSeparator: " "
    shortForm: true
  }
  formatter number #formatterLTR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    emptyValue: "-"
  }
  formatter number #formatterRR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    postfix: " %"
  }

  formatter color #formatterColor {
    thresholds: #009900 >=9 , #b34700 >=7, #b30000 >=0
  }
  formatter color #formatterColor2 {
    thresholds: #0099AA >=9 , #b347AA >=7, #b300AA >=0
  }
  formatter number #metricFormat {
    numberDecimals: 1
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
  }

  formatter number #responsesFormat {
    numberDecimals: 0
    shortForm: false
  }

  formatter color #riskStringFormatter {
    thresholds: Unknown = 0 , Low = 1, Medium = 2, High = 3
  }

  formatter color #valueCases {
    thresholds: #ff0000 >=1, #31363e >=0
  }
  formatter color #backgroundColorFormatter {
    thresholds: #e8f8e0 >= 8.5, #ffeed6 >= 6.5, #fedfe2 >= 0
  }
  formatter color #valueColorFormatter {
    thresholds: #5ba35d >= 8.5, #ffa156 >= 6.5, #dd3435 >= 0
  }
  formatter objectProperty #textPicker {
    property: text
  }

  formatter color #riskColorFormatter {
    thresholds: #FA5263 >= 99%, #FFBD5B >=49%, #82D854 >0%
  }
}

page #AccountList {
  label: "Account List"

  widget markdown {
    size: medium
    markdown: "
## Confirmit Confidential Information"
  }
  widget accountList {
    label: "Accounts"
    table: accounts:
    sortColumn: healthrisk
    sortOrder: descending
    navigateTo: "Account"
    size: large

    hierarchy: accounts:ParentAccountID

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    column hierarchy #accountName {
      label: "Account Name "
      value: accounts:AccountName
      rowHeader: true
    }
    column value #accountMan {
      label: "Account Owner"
      value: accounts:AccountOwner
    }

    column value #healthrisk {
      label: "Health Risk"
      value: IIF(IIF(count(healthCheck:responseid) > 0, 1, 0) = 1, IIF(average(SCORE(healthCheck:Q2)) >= 9, 1, IIF(average(SCORE(healthCheck:Q2)) >= 5, 2, 3)), 0)
      align: center
      format: riskStringFormatter
    }

    column value #relrisk {
      label: "LTR Risk"
      value: IIF(COUNT(respondent:respid) = 0, 0, IIF(IIF(COUNT(survey:responseid, survey:status = "complete" OR survey:status = "incomplete") / COUNT(respondent:respid) * 100 < 5, 0, 1) = 1, IIF(average(SCORE(survey:Q1)) >= 9, 1, IIF(average(SCORE(survey:Q1)) > 6, 2, IIF(average(SCORE(survey:Q1)) > 0, 3, 0))), 0))
      align: center
      format: riskStringFormatter
    }

    column value #revRisk {
      label: "Revenue Risk "
      value: @cp.revenueRiskValue
      align: center
      format: riskStringFormatter
    }

    column metric #hh {
      label: "Health"
      value: average(score(healthCheck:Q2))
      format: formatterLTR
      view: metrics
      target: 9
    }
    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
      align: center
    }

    column value #rev2017 {
      label: "2017 rev"
      value: sum(revenue:AnnualRevenue, revenue:year = 2017)
      format: formatterID
      align: right
    }
    column value #rev2016 {
      label: "2016 rev"
      value: sum(revenue:AnnualRevenue, revenue:year = 2016)
      format: formatterID
      align: right
    }
    column value #revDiff {
      label: "Rev diff"
      value: sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)
      format: formatterID
      align: right
    }
    column value #revDiffPercentage {
      label: "Rev diff"
      value: (sum(revenue:AnnualRevenue, revenue:year = 2017) - sum(revenue:AnnualRevenue, revenue:year = 2016)) / sum(revenue:AnnualRevenue, revenue:year = 2017) * 100
      format: formatterRR
      align: right
    }
    column value #tickets {
      label: "eJournal total"
      value: sum(ejournal:closedTickets)
    }
    column value #ticketsOpen {
      label: "eJournal Open"
      value: sum(ejournal:openTickets)
    }

    column value #case2 {
      label: "Cases"
      value: COUNT(cases:CaseId)
      align: center
      format: responsesFormat

    }
    column value #responses {
      label: "Responses "
      format: valueFMTnses
      value: COUNT(survey:responseid, survey:status = "complete" OR survey:status = "incomplete")
      align: center
    }
    column value #rate {
      label: "Response Rate"
      value: COUNT(survey:responseId, survey:status = "complete" OR survey:status = "incomplete") * 100 / COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
      format: formatterRR
      align: center
    }
    column value #noResp {
      label: "No Response"
      value: COUNT(respondent:respid, respondent:smtpstatus = "messagesent") - COUNT(survey:responseid, survey:status = "Complete")
      align: center
    }
  }
}

page account #Account {
  label: "Account"


  widget search {
    table: accounts:
    layoutArea: "header"
    value: accounts:AccountName + " " + accounts:AccountId
    navigateTo: "AccountPage"
    iconType: "account"
  }

  widget title {
    table: accounts:
    layout column {
      tile value #c {
        value: accounts:accountName
      }
    }
  }

  widget summary {
    size: large
    table: accounts:

    tile metric {
      label: "LTR Average"
      value: average(score(survey:Q1))
      target: 7
    }

    tile metric {
      label: "Health check"
      value: average(score(healthCheck:Q2))
      target: 5
    }


    tile risk {
      label: "Revenue Risk"
        // need to tune formatting! add calculation
      value: @cp.revenueRiskValue
      textValue: IIF(@cp.revenueRiskValue = 3, "High", IIF(@cp.revenueRiskValue = 2, "Medium", IIF(@cp.revenueRiskValue = 1, "Low", "Unknown")))
      min: 1
      max: 3
      target: 0
      renewal: accounts:RenewalDate
      revenue: sum(revenue:AnnualRevenue, revenue:year = 2017)
      backgroundColorFormatter: riskColorFormatter
    }

    tile responseRate {
      invites: COUNT(respondent:respid, respondent:smtpstatus = "messagesent")
      responses: COUNT(survey:responseId, survey:status = "complete" OR survey:status = "incomplete")
    }
  }

  widget contactList #hg {
    size: large
    label: "Contacts "
    table: contacts:
    sortColumn: name
    sortOrder: descending
    navigateTo: "Contact"
    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }
    view metric #ccc {
      valueColorFormatter: valueCases
    }
    column value #name {
      label: "Name"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #company {
      label: "Company"
      value: contacts:AccountName
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }

    column metric #ltr {
      label: "LTR"
      value: average(score(survey:Q1))
      format: formatterLTR
      view: metrics
      target: 9
    }
    column value #openCases {
      label: "Cases"
      value: COUNT(cases:CaseId)
      view: ccc
    }
    column value #lastResponse {
      label: "Last response "
      value: max(survey:interview_start)
      format: date11
      asign: center
    }
    column value #comments {
      label: "Comments"
      value: MAX(survey:Q2, survey:interview_start = max(survey:interview_start))
    }
  }

  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Date"
      value: cases:DateCreated
      align: center
      format: date12
    }

    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000818", "Health Check : At Risk", IIF(cases:Workflow = "1000819", "Health Check : High Potential", "Relationship : Recommend and/or Tech Detractors")))
    }
    column value #res {
      label: "Resolution"
      value: IIF(cases:lk_1548 = "5218" OR cases:lk_1548 = "5219" OR cases:lk_1548 = "5220", "Client specific", IIF(cases:lk_1548 = "5221" OR cases:lk_1548 = "5222" OR cases:lk_1548 = "5223", "Generic", IIF(cases:lk_1548 = "8319" OR cases:lk_1548 = "8320" OR cases:lk_1548 = "8321" OR cases:lk_1548 = "8322", "At risk: Action Taken", IIF(cases:lk_1548 = "8323" OR cases:lk_1548 = "8324", "High potential", "To Be Coded"))))
    }
    column value #link {

      label: "Action"
      value: cases:CaseLink
      view: link1
    }

  }
}

page contact #Contact {
  label: "Contact"


  widget search {
    table: contacts:
    layoutArea: "header"
    value: contacts:client_first_name + " " + contacts:client_last_name
    navigateTo: "Contact"
  }

  widget title {
    table: contacts:
    layout column {
      tile icon {
        value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/magdalenas/defaultLogo.PNG"
      }
    }
    layout column {
      layout row {
        tile value {
          value: contacts:FirstName + " " + contacts:LastName
        }
        tile role {
          value: contacts:ContactRole
        }
      }
      layout row {
        tile company {
          value: contacts:AccountName
        }
      }
    }
  }


  widget summary {
    size: large
    table: contacts:
    tile contactDetails #cc {
      title: contacts:Title
      role: contacts:ContactRole
      email: contacts:email
      phone: contacts:Phone
      industry: contacts:Industry
    }

    tile accountDetails #cc4 {
      accountOwner: contacts:AccountOwner
      salesManager: contacts:SalesLeader1
      region: contacts:WorldRegion
      revenue: contacts:AnnualAccountValue
      renewalDate: accounts:RenewalDate
    }

    tile metric #a {
      label: "LTR"
      value: average(score(survey:Q1))
      target: 7
    }

    tile metric #da {
      label: "Surveys"
      value: count(survey:responseid)
    }
  }

  widget accountCases {
    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Date"
      value: cases:DateCreated
      align: center
      format: date12
    }

    column value #caseSev {
      label: "Status"
      value: IIF(cases:SystemStatus = "Open", "Open", "Closed")
    }
    column value #caseCat {
      label: "Category"
      value: IIF(cases:Workflow = "0", "All attributes and users", IIF(cases:Workflow = "1000818", "Health Check : At Risk", IIF(cases:Workflow = "1000819", "Health Check : High Potential", "Relationship : Recommend and/or Tech Detractors")))
    }
    column value #res {
      label: "Resolution"
      value: IIF(cases:lk_1548 = "5218" OR cases:lk_1548 = "5219" OR cases:lk_1548 = "5220", "Client specific", IIF(cases:lk_1548 = "5221" OR cases:lk_1548 = "5222" OR cases:lk_1548 = "5223", "Generic", IIF(cases:lk_1548 = "8319" OR cases:lk_1548 = "8320" OR cases:lk_1548 = "8321" OR cases:lk_1548 = "8322", "At risk: Action Taken", IIF(cases:lk_1548 = "8323" OR cases:lk_1548 = "8324", "High potential", "To Be Coded"))))
    }
    column value #link {

      label: "CaseLink"
      value: cases:CaseLink
      view: link1
    }

  }
}
title "Sodexo demo"
//Please do not make changes to this report.
//This is a live report shared with the customer

config hub {
  hub: 53071
  table survey = p3080257220.response
  table accounts = crmdata.accounts
  table surveyR = p3080257220.respondent
  table contacts = p3086013448.response
  table acc = crmdata.SHO
  table names = crmdata.ACCNAMES
  relation oneToMany #rel1 {
    primaryKey: accounts:AccountID
    foreignKey: contacts:accountid_crm_formatted
  }
  relation oneToOne #rel2 {
    primaryKey: accounts:district_mgrs
    foreignKey: acc:id
  }
  relation oneToOne #rel3 {
    primaryKey: accounts:AccountID
    foreignKey: names:AccountID
  }
}
config report #cr {
  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Sodexo/Sodexo_logo.jpg"

  formatter number #formatterLTR {
    numberDecimals: 2
    decimalSeparator: "."
  }
  formatter number #formatterRR {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    postfix: "%"
  }
  formatter number #customEmpty {
    numberDecimals: 0
    emptyValue: "-"
  }
  formatter objectProperty #textPicker {
    property: text
  }
  formatter color #backgroundColor {
    thresholds: #e8f8e0 >8, #ffeed6 >6, #fedfe2 >= 0
  }
  formatter color #valueColor {
    thresholds: #388e3c >8, #ff6d00 >6, #d40000 >= 0
  }
  formatter date #DDMMMYYYY {
    format: "DD MMM YYYY"
    shortForm: true
    emptyValue: "-"
  }
  formatter date #dateRelative {
    locale: en
    shortForm: false
    relative: true
  }
  formatter text #commentFormat {
    useDots: true
    length: 68
    emptyValue: "-"
  }
  formatter color #riskSodexo {
    thresholds: #E46C0A >1, #FAC090 > 0, #FFFDFC = 0
  }
  formatter color #riskBgColorFormatter {
    thresholds: #23C813 > 8, #FFAB00 > 6, #ff0000 >= 0
  }
  palette: "#86ABE2","#4079D0","#1B6600","#2D9900","#9CCB00","#FEFE00","#F9BF00","#F18500","#EF6300","#F30000", "#AA0010", "#C0C0C0"

  paletteSod: "#FAC090","#E46C0A"

  formatter number #floatNumber {
    numberDecimals: 1
  }

  formatter date #dateFormat {
    inputFormat: "YYYYMM"
    formatString: "YYYY MMMM"
  }
  formatter text #textDefault1 {
    length: 20
    useDots: true
  }

  state case #currentCase {
    lab: "Case"
    value: COUNT(survey:case_created, survey:case_created = "1")   // AND survey:case_status!='99')
  }
  completeSurv: COUNT(survey:responseid, survey:status = "Complete")
  ltrValue: average(score(survey:Q1.1))
  ltrTarget: 9
  healthTarget: 8
  riskValue: average(SCORE(survey:Q1.1), @cr.currentPeriodFilter)
  riskTarget: 6
  riskSod: IIF(SOME(survey:case_created = "1"), 2, IIF(COUNT(survey:responseid) < 1, 1, 0))
  rateInvites: COUNT(surveyR:respid, surveyR:smtpstatus = "messagesent")
  rateResponses: @cr.completeSurv
  rateValue: @cr.rateResponses / @cr.rateInvites * 100
  casesValue: COUNT(survey:case_created, survey:case_created = "1" AND survey:case_status != "99")
  fullContactName: contacts:client_first_name + " " + contacts:client_last_name
  currentPeriod: max(survey:interview_start) >= 2017-01-01
  previousPeriod: max(survey:interview_start) < 2017-01-01

  currentPeriodFilter: survey:interview_start >= 2017-01-01
  previousPeriodFilter: survey:interview_start < 2017-01-01

}

layoutArea toolbar {
  filter multiselect {
    optionsFrom: survey:survey_method
  }

  filter multiselect {
    optionsFrom: survey:client_contract_role
  }
  filter multiselect {
    optionsFrom: accounts:segment
    label: Segment
  }
  filter multiselect {
    label: "Country"
    optionsFrom: accounts:country
  }
  filter multiselect {
    label: "Region"
    optionsFrom: survey:hRegionCoded
  }
  filter multiselect {
    label: "Account Rating"
    option checkbox {
      label: "Gold"
      value: accounts:revenue > 200000
    }
    option checkbox {
      label: "Silver"
      value: accounts:revenue > 99999 AND accounts:revenue < 199999
    }
    option checkbox {
      label: "Bronze"
      value: accounts:revenue < 100000
    }
  }
  filter multiselect {
    label: "Year"
    option checkbox {
      label: "2017"
      value: survey:interview_start >= 2017-01-01 AND survey:interview_start < 2018-01-01
    }
    option checkbox {
      label: "2016"
      value: survey:interview_start >= 2016-01-01 AND survey:interview_start < 2017-01-01
    }
  }
}

page #Overview {
  label: "Overview"

  widget portfolioBreakdown #z {
    label: "Case Management Risk"
    size: small
    category: Year(survey:interview_start)
    segment: IIF(survey:case_created = "1", "Alert", IIF(IN(survey:status, "incomplete", "notanswered", "quotafull", "error", "screened"), "Silent"))
    value: count(survey:responseid) //, survey:interview_start>2017-01-01)
    palette: @cr.paletteSod

  }
  widget accountList {
    label: "Sites"
    table: accounts:
    size: medium
    sortColumn: case1
    sortOrder: descending
    column value #i {
      label: "Name"
      value: accounts:AccountName
      format: textDefault1
    }
    column value #case1 {
      label: "# of Alerts"
      value: COUNT(survey:case_created, survey:case_created = "1")
      sortable: true
    }
  }
  widget portfolioBreakdown {
    label: "Satisfaction by Segment"
    size: large
    category: survey:segment
    segment: survey:NPS_recode
    value: count(survey:responseId)
    percent: on
  }
  widget portfolioBreakdown #pB {
    label: "Loyalty by month"
    size: large

    category: calendarMonth(survey:interview_start)
    categoryFormat: dateFormat
    value: average(score(survey:Q1.1))
    format: floatNumber
  }

}

page #Sites {
  label: "Sites"

  widget search {
    table: accounts:
    layoutArea: "header"
    value: accounts:AccountName
    navigateTo: Sites

  }
  widget accountList {
    label: "Sites"
    size: large
    table: accounts:
    sortColumn: dd
    sortOrder: descending
    navigateTo: Site
    hierarchy: accounts:HierarchyID
    view icon #icon {
      size: "25"
    }

    column hierarchy #accountName {
      label: "Site"
      value: accounts:AccountName
      rowHeader: true
      format: textDefaultFormatter
    }

    column value #id {
      label: "ID"
      value: accounts:AccountID
    }
    column value #top {
      label: "Top Parent"
      value: accounts:parentid_HierarchyId
    }
    column value #i {
      label: "# Invited (total)"
      value: COUNT(surveyR:respid, surveyR:smtpstatus = "messagesent")
    }
    column value #f {
      label: "# Failed Invites"
      value: COUNT(surveyR:respid, surveyR:smtpstatus = "badmail")
    }
    column value #responses {
      label: "# of Resp"
      value: @cr.completeSurv
    }
    column value #pro {
      label: "# of Promoters"
      value: COUNT(survey:responseid, score(survey:Q1.1) > 8)
    }
    column value {
      label: "# of Passive"
      value: COUNT(survey:responseid, between(score(survey:Q1.1), 7, 8))
    }
    column value #dd {
      label: "# of Detractors"
      value: COUNT(survey:responseid, score(survey:Q1.1) < 7)
    }
    column value {
      label: "# Key Dec Maker Resp"
      value: COUNT(survey:responseid, survey:client_contract_role = "2")

    }
    column value #case1 {
      label: "# of Alerts"
      value: COUNT(survey:case_created, survey:case_created = "1")
      sortable: true
    }
    column value #risk2 {
      label: "Client Loyalty Risk "
      value: IIF(SOME(survey:case_created = "1"), "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/autumnblaze.png", IIF(COUNT(survey:responseid) < 1, "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/sweetorange_r.png", "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Icons%20for%20Studio/transparent.png"))
      view: icon
    }

  }
}


page account #Site {
  label: "Site"

  widget search {
    table: contacts:
    layoutArea: "header"
    value: @cr.fullContactName
    navigateTo: Contact
    hierarchy: accounts:HierarchyID
  }
  widget title {
    table: accounts:
    view camelCSS #subheader {
      color: "rgba(0, 76, 179, 2)"
      marginLeft: "14px"
      fontSize: "18px"
    }
    view camelCSS #subheader2 {
      color: "rgba(13, 24, 33, 0.54)"
      marginLeft: "14px"
      fontSize: "13px"
    }
    layout column {
      tile value {
        value: accounts:AccountName
      }
      tile value {
        value: "VP: " + names:regionvps + "   " + "DM:  " + acc:name
        view: subheader
      }
    }
  }
  widget title #test {
    table: accounts:

    view camelCSS #subheader2 {
      color: "rgba(13, 24, 33, 0.54)"
      marginLeft: "14px"
      fontSize: "13px"
    }
    layout column {
      tile value #c {
        value: "ID: " + accounts:accountId
        view: subheader2
      }
    }
  }

  widget summary {
    table: accounts:
    hierarchy: accounts:HierarchyID

    tile responseRate {
      invites: @cr.rateInvites
      responses: @cr.rateResponses
    }
    tile casesStatus {
      label: "Alerts"
      open: @cr.currentCase.value
      overdue: 0
    }
    tile metric #k {
      label: "Key Dec.Makers"
      value: COUNT(survey:responseid, survey:client_contract_role = "2")
      target: 1

    }
    tile risk {
      label: "Loyalty Risk"
      value: IIF(SOME(survey:case_created = "1"), 2, IIF(COUNT(survey:responseid) < 1, 1, 0))
      target: 1
      min: 0
      max: 2
      renewal: accounts:renewalDate
      revenue: accounts:revenue
      textValue: IIF(SOME(survey:case_created = "1"), "Alert", IIF(COUNT(survey:responseid) < 1, "Silent", " "))
      format: formatterLTR
      backgroundColorFormatter: riskSodexo
    }
  }

  widget contactList {
    label: "Contacts"
    table: contacts:
    inHierarchy: accounts:HierarchyId
    size: large
    sortColumn: company
    sortOrder: ascending
    navigateTo: Contact
    view metricWithChange #metrics {
      backgroundColorFormatter: backgroundColor
      valueColorFormatter: valueColor
      fontSize: small
    }
    column value #name {
      label: "Name"
      value: @cr.fullContactName
    }
    column value #company {
      label: "Site"
      value: accounts:AccountName  //contacts:accountid_crm_formatted
    }

    column metric #ltr {
      label: "Loyalty"
      value: average(score(survey:Q1.1), @cr.currentPeriodFilter)
      previous: average(score(survey:Q1.1), @cr.previousPeriodFilter)
      target: @cr.ltrTarget
      format: formatterLTR
      view: metrics
      align: left
    }

    column value #lastResponse {
      label: "Last Invite Date"
      value: max(survey:InitialInviteDate)
      format: DDMMMYYYY
      align: center
    }
    column value {
      label: "Client Email"
      value: contacts:email

    }

    column value {
      label: "Survey Status"
      value: max(AnswerText(survey:svy_status))

    }

    column value {
      label: "Change\\Resend Status"
      value: max(AnswerText(survey:change_request_status))
    }

    column value #role {
      label: "Role"
      value: contacts:client_contract_role
      format: textPicker
      sortable: false
    }

    column value {
      label: "Alert Status"
      value: max(AnswerText(survey:case_alert_status))
    }
  }
}

page contact #Contact {
  label: "Contact"

  widget search {
    table: accounts:
    layoutArea: "header"
    value: accounts:AccountName + " " + accounts:accountid_crm_formatted
    navigateTo: Account
    iconType: "account"
  }
  widget title {
    table: contacts:
    view icon #ii {
      size: "65"
      roundedCorner: true

    }
    layout column {
      tile value #firstName {
        value: contacts:client_first_name
      }
      tile value #lastName {
        value: contacts:client_last_name
      }
      tile value #role {
        value: contacts:client_contract_role
        format: textPicker
      }
      tile value #account {
        value: accounts:AccountName
      }
      tile icon {
        value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Confirmit%20new%20layout/53633418-5037-4CEB-AF68-D8616D95094B.jpg"
        view: ii
      }
    }
  }
  widget summary {
    size: large
    table: contacts:
    tile contactDetails #cc {
      email: contacts:email
      title: contacts:contact_title
      phone: contacts:client_phone
      role: AnswerText(contacts:client_contract_role)
      industry: max(AnswerText(accounts:segment))
    }
    tile accountDetails #cc4 {
      accountOwner: names:regionvps //(accounts:area_vps + " (") + (accounts:alert_email + ")")
      salesManager: names:districtmgrs
      region: max(survey:region)
      revenue: accounts:revenue
      renewalDate: accounts:RenewalDate
    }
    tile metric {
      label: "LTR"
      value: average(score(survey:Q1.1))
      target: 9
    }
    tile surveyResponses #da {
      label: "Survey Responses"
      total: count(survey:responseid)
      completed: @cr.completeSurv
    }
    tile casesStatus {
      open: COUNT(survey:case_created, survey:case_created = "1")
      overdue: 0
    }
  }
  widget contactSurveys {
    label: "Surveys"
    table: survey:
    view metricWithChange #metrics {
      backgroundColorFormatter: backgroundColor
      valueColorFormatter: valueColor
      fontSize: small
    }
    sortColumn: s6
    size: large
    sortOrder: ascending


    column value #s2 {
      label: "Status"
      value: survey:status
    }

    column value #is {
      label: "Date"
      value: survey:interview_start
      format: DDMMMYYYY
    }

    column metric #s3 {
      label: "LTR"
      value: average(score(survey:Q1.1), @cr.currentPeriodFilter)
      previous: average(score(survey:Q1.1), @cr.previousPeriodFilter)
      target: @cr.ltrTarget
      format: formatterLTR
      align: center
      view: metrics

    }

    column value #cc {
      label: "Cases"
      value: @currentCase.value

    }
    column value #s5 {
      label: "email"
      value: survey:email
    }

    column value #s6 {
      label: "comments"
      value: survey:Q8
      format: commentFormat
    }

  }

  widget accountCases {
    label: "Cases"
    table: survey:
    size: large
    sortColumn: caseid
    sortOrder: ascending
    column value #lastResponse {
      label: "Date"
      value: survey:ResponseEndDate
      format: DDMMMYYYY
    }
    column value #caseid {
      label: "Cases"
      value: COUNT(survey:case_created, survey:case_created = "1")
    }

    column value #cas {
      label: "Status"
      value: survey:case_status
      format: textPicker
    }
    column value #alert {
      label: "Alert"
      value: survey:case_alert_status
      format: textPicker
    }
    column value #caseSev {
      label: "Case Status Final"
      value: survey:case_status_final
      format: textPicker
    }
  }
}



state url #urlParams {
  surveyResponseTable: ""
}

config hub {
  hub: 123
  table survey = @urlParams.surveyResponseTable

  dimensionGroup #favNeuNonFav {

    dimension #engagement {
      label: "Engagement"
      questions: s1, s2, s3, s4, s5NotRequired, m1, m2
    }

    dimension #ethicsAndCompliance {
      label: "Ethics & Compliance"
      questions: s6, s7, s8, s9
    }

    dimension #safety {
      label: "Safety"
      questions: s10, s11, s12, s13
    }

    dimension #openness {
      label: "Openness"
      questions: i1, i2LongText, t1, t2NotRequired, t3LongText, s14LongText
    }

    option favorable {
      label: "Favorable"
      score: 100
    }

    option neutral {
      label: "Neutral"
      score: 50
    }
    option nonFavorable {
      label: "Non-favorable"
      score: 0
    }

    recodingRule #fivePoint {
      mapping {
        to: favorable
        from: 1,2
      }
      mapping {
        to: neutral
        from: 3
      }
      mapping {
        to: nonFavorable
        from: 4,5
      }
    }

    recodingRule #fivePointFlipped {
      mapping {
        to: favorable
        from: 4,5
      }
      mapping {
        to: neutral
        from: 3
      }
      mapping {
        to: nonFavorable
        from: 1,2
      }
      questions: s5NotRequired, s6
    }

    defaultRecodingRule: fivePoint
  }

  dimensionGroup #WPA {
    dimension #WPA {
      label: "WPA"
      questions: s50, m52
    }
  }
}

config pulse {
  workflowPage: "workflow"
  overviewPage: "overview"
  reportPage: "report"
  wpaPage: "wpa"
  surveyListPage: "surveylist"
  reportAccessPage: "reportaccess"

  librarySurvey: p1230235
  contactDatabase: p1230087
  languages: en, no

  minNumberOfRecipients: 10
  maxNumberOfRecipients: 60

  surveyDurationInDays: 9
  sendInSelectedLanguageOnly: false
  delayDaysBeforeFirstReminder: 2
  delayDaysBeforeSubsequentReminders: 2
  totalReminders: 3
  minutesBetweenBatches: 30
  batchSize: 100

  dimensionStyle {
    dimension: engagement
    description: "Describe the category here"
    color: green
    icon: "rowing"
  }

  dimensionStyle {
    dimension: ethicsAndCompliance
    description: "Describe the category here"
    color: blue
    icon: "office-building"
  }

  dimensionStyle {
    dimension: safety
    description: "Describe the category here"
    color: blue
    icon: "hearing"
  }

  dimensionStyle {
    dimension: openness
    description: "Describe the category here"
    color: blue
    icon: "bubble_chart"
  }

  dimensionStyle {
    dimension: WPA
    description: "Describe the category here"
    color: blue
    icon: "bubble_chart"
  }

  template pulse #ecd {
    label: "Engagement & Career Development"
    notes: "This survey focuses on employees' commitment and advocacy for the company as a place to work and their insights into future development at the company."
    locked: true
    questions: s1, s2, s3, s4, s5NotRequired, m1, m2
    lockedQuestions: s1, s2, s3, s4, s5NotRequired, m1, m2
    languages: en, no
    emailInvite: e1
    emailReminder: e2
  }

  template pulse #organizationalCulture {
    label: "Organizational Culture"
    notes: "These questions measure perceptions of quality of products and services, commitment to delivering high quality products and services and innovation of products."
    questions: s6, s7, s8, s9
    lockedQuestions: s6
    languages: en
    emailInvite: e1
  }

  template pulse #safety {
    label: "Safety"
    notes: "These questions measure perceptions of safety at work."
    questions: s10, s11, s12
    emailInvite: e1
  }

  template pulse #openness {
    label: "Openness"
    notes: "These questions measure perceptions of openness at work."
    questions: i1, i2LongText, t1, t2NotRequired, t3LongText, s14LongText
    emailInvite: e1
  }

  template pulse #WPA {
    label: "Work Place Assessment"
    notes: "Work Place Assessment."
    locked: true
    questions: s50, m52
    lockedQuestions: s50, s52
    languages: en
    emailInvite: e1
    emailReminder: e2
  }
}

config sampling {
  filter hierarchy {
    question: hierarchy
  }

  filter multiselect {
    question: location
  }
}

page #workflow {
  label: "workflow"

  hide: true
  widget workflowHeader {
    layoutArea: "header"
  }

  widget agileWorkflow {
    label: "Workflow"

    step reviewTemplate #Reviewtemplate

    step customize #Customize

    step selectSample #Selectsample {
      widget sampling {

      }
    }

    step setUpEmail #Setupemail {

    }

    step commit #Commit {
      widget samplingInfo
    }
  }
}

page #surveylist {
  label: "Surveys"

  widget agileHeader {
    layoutArea: "header"
  }

  widget surveyList {
    name: "testname"
    label: "Survey list"
  }
}

page #library {
  label: "Survey Library"

  widget agileHeader {
    layoutArea: "header"
  }

  widget templateList
}


page #overview {
  hide: true
  label: "Survey Overview"

  widget agileHeader {
    layoutArea: "header"
    hideNewSurvey: true
    showBackButton: true
  }

  widget surveyOverview {
    widget responseOverview {

    }

    widget surveyCalendar {

    }
  }
}

page #report {
  hide: true
  label: "Survey Report"

  widget agileHeader {
    layoutArea: "header"
    hideNewSurvey: true
    showBackButton: true
  }

  widget surveyReport {
    widget responseOverview {

    }

    widget surveyScores {
      dimensionGroup: favNeuNonFav
    }

    widget surveyComments {

    }
  }
}

page #reportaccess {
  hide: true
  label: "Sharing"

  widget agileHeader {
    layoutArea: "header"
    hideNewSurvey: true
    showBackButton: true
  }

  widget reportAccess {
  }
}


page #wpa {
  hide: true
  label: "Work Place Assessment"
  widget agileHeader {
    layoutArea: "header"
  }


  widget questionBreakdown {
    label: "Violence, threats, bullying and harassment"
    percent: on
    question: survey:m52
    mode: barchart
  }

  widget questionsScores {
    view itemBar #questionsScoresItemBarDefaultView
    label: "Psychosocial working environment"
    size: large
    tile list {
      item bar { question: survey:s50 }
    }
  }
}

config access {
  portalid: 123
}