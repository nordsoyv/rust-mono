title "Frank Empower test"


// //APPLY SSO FROM SALESFORCE
// config access {
//   portalid: 1870
//   ssoConfig: Confirmit_Salesforce
// }

config editor {
  trace: true
}

config queryOptions {
  optimization {
    CachingProfitLimit: "0"
  }
}

//CONFIGURE HUB
config hub {
  hub: 4203
  numRequests: 3
//FEEDBACK SOURCES
  table relationship = relationship.response  //relationship survey
  table respondent = relationship.respondent  //relationship respondent
  table teamcheck = teamcheck.response  //internal team check survey
  table teamcheckresp = teamcheck.respondent //internal team check respondent
  table website = website.response //www.confirmit.com feedback survey
  table clientandteam = combinedREL_TC.response //relationpgeship + teamcheck combined

  table feedback = p1879470485.response // EMPOWER feedback survey

  //CONTACT DB
  table contacts = contacts.response // contact database

  //FINANCE£
  table finance = EmpowerKPI.EmpowerKPI //Internal finance team results

  //EJOURNAL DATA
  table TicketSummary = eJournal.TicketSummary
  table TicketCategories = eJournal.TicketCategories

  //SFDC
  table SFDCAccounts = fromcrmconnector.SFDCAccounts_v6_0_1
  table SFDCHorizonsSites = fromcrmconnector.SFDCHorizonsSites_v6_0_1
  table SFDCMarketLeads = fromcrmconnector.SFDCContactMktoLeadScore
  table SFDCClosedOpportunities = fromcrmconnector.FiveYrsClosedOpportunities_v6_0_1
  table SFDCeJournalAccounts = fromcrmconnector.SFDCeJournalAccounts_v6_0_1

  //HORISONS ACCOUNT OVERVIEW DATA
  table usageAccounts = crmdata_combined.Accounts
  table usageAccountStatistics = crmdata_combined.AccountStatistics
  table usageActivatedModules = crmdata_combined.ActivatedModules
  table usageFlexExtensions = crmdata_combined.FlexExtensions
  table usageLicenses = crmdata_combined.Licenses
  table usageProfessionalUsers = crmdata_combined.ProfessionalUsers
  table usageReportalLicenses = crmdata_combined.ReportalLicenses
  table usageStandardUsers = crmdata_combined.StandardUsers
  table usageTranslatorUsers = crmdata_combined.TranslatorUsers


  //ACTIONs
  table cases = am.CASE //ACTION MANAGEMENT
  table apInitiatives = ap.initiative //ACTION PLANNER

  //HIERARCHIES
  table hierarchy = dbdesigner.21039

  //hierarchy --> accounts
  relation oneToMany {
    primaryKey: hierarchy:id
    foreignKey: SFDCAccounts:id
  }

  // accounts --> Team Check respondent --> Team Check Survey
  relation oneToMany {
    primaryKey: SFDCAccounts:id
    foreignKey: teamcheckresp:AccountID
  }

  // accounts --> contact db
  relation oneToMany {
    primaryKey: SFDCAccounts:id
    foreignKey: contacts:AccountID
  }
  //accounts to market leads
  relation oneToMany {
    primaryKey: SFDCAccounts:id
    foreignKey: SFDCMarketLeads:AccountId
  }

  //eJOURNAL ACCOUNT RELATIONSHIPS
  relation oneToMany #relSFDCeJournalAccounts {
    primaryKey: SFDCAccounts:Id
    foreignKey: SFDCeJournalAccounts:AccountID
  }
  relation oneToMany #eJournalTicketSummary {
    primaryKey: SFDCeJournalAccounts:eJournalAccountID
    foreignKey: TicketSummary:CompanyId
  }
  relation oneToMany #eJournalTicketCategory {
    primaryKey: TicketSummary:CategoryId
    foreignKey: TicketCategories:id
  }

  //HORISONS ACCOUNT OVERVIEW RELATIONSHIPS
  relation oneToMany #relSFDCHorizonsSites {
    primaryKey: SFDCAccounts:Id
    foreignKey: SFDCHorizonsSites:AccountID
  }

  relation oneToMany #relSFDCClosedOpportunities {
    primaryKey: SFDCAccounts:Id
    foreignKey: SFDCClosedOpportunities:AccountId
  }

  relation oneToMany #relHorizonsSitesToUsageAccounts {
    primaryKey: SFDCHorizonsSites:CompositeAccountID
    foreignKey: usageAccounts:CompositeAccountId
  }

  relation oneToMany #relUsageAccountStatistics {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageAccountStatistics:CompositeAccountId
  }

  relation oneToMany #relUsageActivatedModules {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageActivatedModules:CompositeAccountId
  }

  relation oneToMany #relUsageFlexExtentions {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageFlexExtensions:CompositeAccountId
  }

  relation oneToMany #relUsageLicenses {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageLicenses:CompositeAccountId
  }

  relation oneToMany #relUsageProfessionalUsers {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageProfessionalUsers:CompositeAccountId
  }

  relation oneToMany #relUsageReportalLicenses {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageReportalLicenses:CompositeAccountId
  }

  relation oneToMany #relUsageStandardUsers {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageStandardUsers:CompositeAccountId
  }

  relation oneToMany #relUsageTranslatorUsers {
    primaryKey: usageAccounts:CompositeAccountId
    foreignKey: usageTranslatorUsers:CompositeAccountId
  }

  //DERIVED VARIABLES
  //For response rate reporting
  variable singleChoice #responseStatus {
    table: respondent:
    label: "Status"
    value: IIF(@filter.isResponded, "c", IIF(@filter.isOptOut, "o", IIF(@filter.isPartial, "p", IIF(@filter.isFailedInvite, "f", "n"))))

    option code {
      code: "f"
      label: "Failed invites"
    }

    option code {
      code: "o"
      label: "Opt-Outs"
    }

    option code {
      code: "n"
      label: "Not responded"
    }

    option code {
      code: "p"
      label: "Partial response"
    }

    option code {
      code: "c"
      label: "Full response"
    }

  }

  variable singleChoice #overdue {
    label: "Overdue"
    table: cases:
    value: IIF(cases:DateDue < GetDate(), "Overdue", "Not")

    option code {
      code: "not"
      score: 1
      label: "No"
    }
    option code {
      code: "overdue"
      score: 2
      label: "Yes"
    }
  }


  variable singleChoice #sClientType {
    label: "Client Type"
    table: SFDCAccounts:
    option code {
      code: "MR"
      score: 1
      label: "MR"
    }
    option code {
      code: "VoC"
      score: 2
      label: "VoC"
    }
    option code {
      code: "VoE"
      score: 3
      label: "VoE"
    }
    option code {
      code: "Unknown"
      score: 4
      label: "Unknown"
    }
    value: IIF(SFDCAccounts:ClientType = "MR", "MR", IIF(SFDCAccounts:ClientType = "VoC", "VoC", IIF(SFDCAccounts:ClientType = "VoE", "VoE", "Unknown")))
  }

  variable singleChoice #sTypeOfCustomer {
    label: "Type of Customer"
    table: SFDCAccounts:
    option code {
      code: "1"
      score: 1
      label: "Self service"
    }
    option code {
      code: "2"
      score: 2
      label: "Hybrid"
    }
    option code {
      code: "3"
      score: 3
      label: "Managed Services"
    }
    option code {
      code: "4"
      score: 4
      label: "Panel / Sample provider"
    }

    option code {
      code: "5"
      score: 5
      label: "Fieldwork agency"
    }

    option code {
      code: "6"
      score: 6
      label: "Full Service Agency"
    }

    option code {
      code: "7"
      score: 7
      label: "Outsourcing / Scripting Services"
    }

    option code {
      code: "Unknown"
      score: 7
      label: "Unknown"
    }

    value: IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "1", "1", IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "2", "2", IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "3", "3", IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "4", "4", IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "5", "5", IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "6", "6", IIF(Last(teamcheck:Q13, teamcheck:interview_start) = "7", "7", "Unknown")))))))
  }

  variable singleChoice #sAccountTeam {
    label: "Account Team"
    table: SFDCAccounts:
    option code {
      code: "1"
      score: 1
      label: "1) Nordic VoC"
    }
    option code {
      code: "2"
      score: 2
      label: "2) EMEA VoC"
    }
    option code {
      code: "3"
      score: 3
      label: "3) EMEA MR"
    }
    option code {
      code: "4"
      score: 4
      label: "4) Russia"
    }

    option code {
      code: "5"
      score: 5
      label: "5) APAC"
    }

    option code {
      code: "6"
      score: 6
      label: "6) US VoC"
    }

    option code {
      code: "7"
      score: 7
      label: "7) Global VoE"
    }

    option code {
      code: "8"
      score: 8
      label: "8) US MR"
    }

    option code {
      code: "Unkown"
      score: 9
      label: "Unkown"
    }
    value: IIF(SFDCAccounts:SalesRegion = "1) Nordic VoC", "1", IIF(SFDCAccounts:SalesRegion = "2) EMEA VoC", "2", IIF(SFDCAccounts:SalesRegion = "3) EMEA MR", "3", IIF(SFDCAccounts:SalesRegion = "4) Russia", "4", IIF(SFDCAccounts:SalesRegion = "5) APAC", "5", IIF(SFDCAccounts:SalesRegion = "6) US VoC", "6", IIF(SFDCAccounts:SalesRegion = "7) Global VoE", "7", IIF(SFDCAccounts:SalesRegion = "8) US MR", "8", "Unknown"))))))))
  }

    //DERIVED VARIABLES
  // variable auto #currActiveUser {
  //   table: SFDCAccounts:
  //   value: sum(usage:uniqueLogins, InMonth(usage:Month, -1, -1))
  //   label: "Current Active Users"
  // }
  // variable auto #prevActiveUser {
  //   table: SFDCAccounts:
  //   value: sum(usage:uniqueLogins, InMonth(usage:Month, -2, -2))
  //   label: "Previous Active Users"
  // }

  variable auto #LastRespondentId {
    table: contacts:
    value: Last(respondent:respid, respondent:FirstEmailedDate, respondent:ContactID = contacts:ContactID)
  }
  variable auto #usersLicenses {
    table: SFDCAccounts:
    value: sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)")
    label: "Users - Licenses"
  }
  variable auto #usersAssigned {
    table: SFDCAccounts:
    value: sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)")
    label: "Users - Assigned"
  }
  variable auto #usages {
    table: SFDCAccounts:
    value: round(IIF(SFDCAccounts:usersLicenses > 0, SFDCAccounts:usersAssigned / SFDCAccounts:usersLicenses * 100), 1)
    label: "Usages"
  }
  variable auto #respCount {
    table: SFDCAccounts:
    label: "Respondent Count"
    value: COUNT(respondent:respid)
  }
  variable auto #FutureBCCCP {
    table: SFDCAccounts:
    value: Sum(SFDCClosedOpportunities:Amount_USD, SFDCClosedOpportunities:CloseDate > GetDate())
    label: "Best Case / Closed / Commit / Pipeline"
  }
  variable auto #ltrL12MRev {
    table: SFDCAccounts:
    value: Sum(SFDCClosedOpportunities:Amount_USD, Between(SFDCClosedOpportunities:CloseDate, AddYear(GetDate(), -1), GetDate()) AND SFDCClosedOpportunities:IsClosed = "true")
    label: "Last 12 mths Revenue"
  }
  variable auto #ltrP12MRev {
    table: SFDCAccounts:
    value: Sum(SFDCClosedOpportunities:Amount_USD, Between(SFDCClosedOpportunities:CloseDate, AddYear(GetDate(), -2), AddYear(GetDate(), -1)) AND SFDCClosedOpportunities:IsClosed = "true")
    label: "Previous 12 mths Revenue"
  }
  variable auto #revDiff {
    table: SFDCAccounts:
    value: round((SFDCAccounts:ltrL12MRev - SFDCAccounts:ltrP12MRev) / SFDCAccounts:ltrL12MRev * 100, 2)
    label: "Revenue Difference"
  }
  variable auto #responseRateL12M {
    table: SFDCAccounts:
    value: round(COUNT(relationship:responseId, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRelRate) * 100 / COUNT(respondent:respid, @filter.isSent AND @daterange.L12MonthRelResp), 1)
    label: "Last 12 mths Response Rate"
  }
  variable auto #noResponsesL12M {
    table: SFDCAccounts:
    value: COUNT(relationship:responseId, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRelRate)
    label: "Last 12 mths no Responses"
  }
  variable auto #invitedL12M {
    table: SFDCAccounts:
    value: COUNT(respondent:respid, @filter.isSent AND @daterange.L12MonthRelResp)
    label: "Invited in Last 12 mths"
  }
  variable auto #NPSavg {
    table: SFDCAccounts:
    value: round(average(score(relationship:Q1), @daterange.L12MonthRel), 1)
    label: "NPS average in Last 12 mths"
  }
  variable auto #NEEDSavg {
    table: SFDCAccounts:
    value: round(average(score(relationship:Q12), @daterange.L12MonthRel), 1)
    label: "Needs average in Last 12 mths"
  }
  variable auto #VALUEavg {
    table: SFDCAccounts:
    value: round(average(score(relationship:Q3), @daterange.L12MonthRel), 1)
    label: "Value average in Last 12 mths"
  }
  variable auto #RELavg {
    table: SFDCAccounts:
    value: round(average(score(relationship:Q4), @daterange.L12MonthRel), 1)
    label: "Relationship average in Last 12 mths"
  }
  variable auto #TECHavg {
    table: SFDCAccounts:
    value: round(average(score(relationship:Q7), @daterange.L12MonthRel), 1)
    label: "Technology average in Last 12 mths"
  }
  variable auto #tNPSavg {
    table: SFDCAccounts:
    value: last(score(teamcheck:Q1), teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC)
    label: "Team NPS average in Last 12 mths"
  }
  variable auto #RENEWavg {
    table: SFDCAccounts:
    value: last(score(teamcheck:Q2), teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC)
    label: "Renew average in Last 12 mths"
  }
  variable auto #BENavg {
    table: SFDCAccounts:
    value: last(score(teamcheck:Q8), teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC)
    label: "Benefits average in Last 12 mths"
  }
  variable auto #EXPavg {
    table: SFDCAccounts:
    value: last(score(teamcheck:Q9), teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC)
    label: "Experience average in Last 12 mths"
  }
  variable auto #sumOfClientWeight {
    table: SFDCAccounts:
    value: IIF(SFDCAccounts:NPSavg >= 0, @weight.NPS, 0) + IIF(SFDCAccounts:NEEDSavg >= 0, @weight.Needs, 0) + IIF(SFDCAccounts:VALUEavg >= 0, @weight.Value, 0) + IIF(SFDCAccounts:RELavg >= 0, @weight.Relationship, 0) + IIF(SFDCAccounts:TECHavg >= 0, @weight.Technology, 0)
    label: "Sum of Client Feeling Weights"
  }
  variable auto #clientFeelingIndex {
    table: SFDCAccounts:
    value: round(IIF(SFDCAccounts:sumOfClientWeight > 0, (IIF(SFDCAccounts:NPSavg >= 0, @index.NPS * @weight.NPS, 0) + IIF(SFDCAccounts:NEEDSavg >= 0, @index.Needs * @weight.Needs, 0) + IIF(SFDCAccounts:VALUEavg >= 0, @index.Value * @weight.Value, 0) + IIF(SFDCAccounts:RELavg >= 0, @index.Relationship * @weight.Relationship, 0) + IIF(SFDCAccounts:TECHavg >= 0, @index.Technology * @weight.Technology, 0)) / SFDCAccounts:sumOfClientWeight), 1)
    label: "Client Feeling Index"
  }

  variable auto #clientFeelingRiskCategory {
    table: SFDCAccounts:
    value: IIF(SFDCAccounts:clientFeelingIndex >= 0, IIF(SFDCAccounts:clientFeelingIndex >= 9, "Low", IIF(SFDCAccounts:clientFeelingIndex >= 7, "Med", "High")), "Unknown")
    label: "Client Feeling Risk Category"
  }

  variable auto #sumOfTeamWeight {
    table: SFDCAccounts:
    value: IIF(SFDCAccounts:tNPSavg >= 0, @weight.tNPS, 0) + IIF(SFDCAccounts:RENEWavg >= 0, @weight.Renew, 0) + IIF(SFDCAccounts:BENavg >= 0, @weight.Benefits, 0) + IIF(SFDCAccounts:EXPavg >= 0, @weight.Experience, 0)
    label: "Sum of Team Feeling Weights"
  }
  variable auto #teamFeelingIndex {
    table: SFDCAccounts:
    value: round(IIF(SFDCAccounts:sumOfTeamWeight > 0, (IIF(SFDCAccounts:tNPSavg >= 0, @index.tNPS * @weight.tNPS, 0) + IIF(SFDCAccounts:RENEWavg >= 0, @index.Renew * @weight.Renew, 0) + IIF(SFDCAccounts:BENavg >= 0, @index.Benefits * @weight.Benefits, 0) + IIF(SFDCAccounts:EXPavg >= 0, @index.Experience * @weight.Experience, 0)) / SFDCAccounts:sumOfTeamWeight), 1)
    label: "Team Feeling Index"
  }

  variable auto #teamFeelingRiskCategory {
    table: SFDCAccounts:
    value: IIF(SFDCAccounts:teamFeelingIndex >= 0, IIF(SFDCAccounts:teamFeelingIndex >= 9, "Low", IIF(SFDCAccounts:teamFeelingIndex >= 7, "Med", "High")), "Unknown")
    label: "Team Feeling Risk Category"
  }

  variable auto #sumOfBehaviourWeight {
    table: SFDCAccounts:
    value: IIF(@index.SpendTrend >= 0, @weight.SpendTrend, 0) + IIF(@index.UserAdoption >= 0, @weight.UserAdoption, 0) + IIF(@index.LeadScore >= 0, @weight.LeadScore, 0) + IIF(@index.ResponseRate >= 0, @weight.ResponseRate, 0)
    label: "Sum of Client Behaviour Weights"
  }
  variable auto #clientBehaviourIndex {
    table: SFDCAccounts:
    value: round(IIF(SFDCAccounts:sumOfBehaviourWeight > 0, (IIF(@index.ResponseRate >= 0, @index.ResponseRate * @weight.ResponseRate, 0) + IIF(@index.SpendTrend >= 0, @index.SpendTrend * @weight.SpendTrend, 0) + IIF(@index.LeadScore >= 0, @index.LeadScore * @weight.LeadScore, 0) + IIF(@index.UserAdoption >= 0, @index.UserAdoption * @weight.UserAdoption, 0)) / SFDCAccounts:sumOfBehaviourWeight), 1)
    label: "Client Behaviour Index"
  }

  variable auto #clientBehaviourRiskCategory {
    table: SFDCAccounts:
    value: IIF(SFDCAccounts:clientBehaviourIndex >= 0, IIF(SFDCAccounts:clientBehaviourIndex >= 9, "Low", IIF(SFDCAccounts:clientBehaviourIndex >= 7, "Med", "High")), "Unknown")
    label: "Client Behaviour Risk Category"
  }
  variable auto #sumOfOverallWeight {
    table: SFDCAccounts:
    value: IIF(SFDCAccounts:clientFeelingIndex >= 0, @weight.clientfeeling, 0) + IIF(SFDCAccounts:teamFeelingIndex >= 0, @weight.teamfeeling, 0) + IIF(SFDCAccounts:clientBehaviourIndex >= 0, @weight.doing, 0)
    label: "Sum of Team Overall Weights"
  }
  variable auto #overallIndex {
    table: SFDCAccounts:
    value: round(IIF(SFDCAccounts:sumOfOverallWeight > 0, (IIF(SFDCAccounts:clientFeelingIndex >= 0, SFDCAccounts:clientFeelingIndex * @weight.clientfeeling, 0) + IIF(SFDCAccounts:teamFeelingIndex >= 0, SFDCAccounts:teamFeelingIndex * @weight.teamfeeling, 0) + IIF(SFDCAccounts:clientBehaviourIndex >= 0, SFDCAccounts:clientBehaviourIndex * @weight.doing, 0)) / SFDCAccounts:sumOfOverallWeight), 1)
    label: "Overall Index"
  }
  variable auto #overallHealthRiskCategory {
    table: SFDCAccounts:
    value: IIF((SFDCAccounts:clientFeelingRiskCategory = "High" AND SFDCAccounts:clientBehaviourRiskCategory = "High") AND (SFDCAccounts:teamFeelingRiskCategory = "High" OR SFDCAccounts:teamFeelingRiskCategory = "Unknown"), "Priority 1", IIF(_IsNull(SFDCAccounts:overallIndex), "Unknown", IIF(SFDCAccounts:overallIndex >= 8, "Priority 4", IIF(SFDCAccounts:overallIndex >= 6, "Priority 3", "Priority 2"))))
    label: "Overall Health Risk Category"
  }

// NOT IN USE AT THE MOMENT (SIMPLIFIED MODEL)
  // variable auto #sumOfOverallWeight2 {
  //   table: accounts:
  //   value: IIF(accounts:clientFeelingIndex >= 0, @weight.clientfeeling2, 0) + IIF(accounts:teamFeelingIndex >= 0, @weight.teamfeeling2, 0)
  //   label: "Sum of Team Overall Weights (simplified)"
  // }
  // variable auto #overallIndex2 {
  //   table: accounts:
  //   value: IIF(accounts:sumOfOverallWeight2 > 0, (IIF(accounts:clientFeelingIndex >= 0, accounts:clientFeelingIndex * @weight.clientfeeling2, 0) + IIF(accounts:teamFeelingIndex >= 0, accounts:teamFeelingIndex * @weight.teamfeeling2, 0)) / accounts:sumOfOverallWeight2)
  //   label: "Overall Index (simplified)"
  // }
  // variable auto #overallHealthRiskCategory2 {
  //   table: accounts:
  //   value: IIF(accounts:teamFeelingRiskCategory = "High" AND (accounts:teamFeelingRiskCategory = "High" OR accounts:teamFeelingRiskCategory = "Unknown"), "High Risk", IIF(_IsNull(accounts:overallIndex2), "Unknown", IIF(accounts:overallIndex2 >= 8, "Secure", IIF(accounts:overallIndex2 >= 6, "Low Risk", "Vulnerable"))))
  //   label: "Overall Health Risk Category (simplified)"
  // }

  variable singleChoice #accountActivityStatus {
    label: "Active and/or Surveyed"
    table: SFDCAccounts:

    option code {
      code: "1"
      score: 1
      label: "Active and/or Surveyed"
    }
    option code {
      code: "2"
      score: 2
      label: "InActive and not surveyed"
    }
    value: IIF((COUNT(respondent:respid, @daterange.L12MonthRelResp AND @filter.isSent) > 0 OR COUNT(teamcheckresp:respid, @daterange.L12MonthTCResp AND @filter.isTeamSent) > 0) OR SFDCAccounts:ActiveClient = "True", "1", "2")
  }

  variable singleChoice #riskgroups {
    label: "Risk"
    table: SFDCAccounts:
    option code {
      code: "Priority 1"
      score: 4
      label: "Priority 1"
    }
    option code {
      code: "Priority 2"
      score: 3
      label: "Priority 2"
    }
    option code {
      code: "Priority 3"
      score: 2
      label: "Priority 3"
    }
    option code {
      code: "Priority 4"
      score: 1
      label: "Priority 4"
    }
    option code {
      code: "Unknown"
      score: 0
      label: "Unknown"
    }
    value: SFDCAccounts:overallHealthRiskCategory

  }
}
//END CONFIGURE HUB SOURCES FOR USE IN THIS REPORT****************************************************************************************

drillDown #accountOwner {

  filter expression {
    value: IIF(SFDCAccounts:accountActivityStatus = "1", true, false)
  }
  level distinct {
    table: SFDCAccounts:
    value: SFDCAccounts:AccountOwnerName
  }
}

drillDown #salesRegion {
  level distinct {
    table: SFDCAccounts:
    value: SFDCAccounts:SalesRegion
  }
}

//REPORT PROPERTIES
config report {

  logo: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/EMPOWER/EmpowerLogo_dk.png"

  //NUMERIC & DATE FORMATS
  formatter date #long {
    formatString: "DD MMM YYYY"
    emptyValue: "None"
  }
  formatter date #monthlabel {
    inputFormat: "YYYYMM"
    formatString: "MMM 'YY"
  }

  formatter date #quarterlabel {
    inputFormat: "YYYYQQ"
    formatString: "'YY Qo"
  }

  formatter value #emptyvalue {
    emptyValue: " "
  }
  formatter number #UScurrency {
    numberDecimals: 0
    prefix: "$ "
    //decimalSeparator: ""
    integerSeparator: ","
    shortForm: true
  }
  formatter number #nodecimal {
    numberDecimals: 0
    decimalSeparator: ""
    integerSeparator: ","
    //shortForm: true
    emptyValue: "-"
  }

  formatter number #nodecimalblank {
    numberDecimals: 0
    decimalSeparator: "."
    shortForm: true
    emptyValue: "NA"
  }

  formatter number #onedecimal {
    numberDecimals: 1
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
  }
  formatter number #twodecimal {
    numberDecimals: 2
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
  }

  formatter number #percentage {
    numberDecimals: 0
    decimalSeparator: "."
    postfix: " %"
  }
  formatter number #percentageonedecimal {
    numberDecimals: 1
    decimalSeparator: "."
    postfix: " %"
  }

  //STYLES: COLOR PALETTES & CONDITIONAL FORMATTING

  //COLOR PALETTES
  formatter color #metricbar {
    thresholds: #0F5E7D >= 1
  }

  //CONDITIONAL FORMATTING
  formatter color #npsGauge {
    thresholds: #82D854 >= 20, #FFBD5B >= 10, #FA5263 >=-100
  }
  formatter color #NetSalesGauge {
    thresholds: #82D854 >= 100, #FFBD5B >= 95,#FA5263 >= 0
  }
  formatter color #RenewalRateGauge {
    thresholds: #82D854 >= 95, #FFBD5B >= 90,#FA5263 >= 0
  }
  formatter color #acrossTheJourney {
    thresholds: #82D854 >= 8, #ffa156 >= 6.5, #dd3435 >= 0
  }
  formatter color #riskleveltextcolor {
    thresholds: #FFFFFF >=9, #333333 >=5, #FFFFFF <5
  }
  formatter color #backgroundColorFormatter {
    thresholds: rgba(126, 210, 81, 0.655) >=9, rgba(255, 187, 92, 0.765) >= 7, rgba(247, 99, 114, 0.731) >= 0
  }
  formatter color #backgroundColorFormatterIndex {
    thresholds: #7ED251 >=8, #FFBB5C >= 6, #F76373 >= 0,#E0E0E0 <0
    defaultValue: transparent
  }
  formatter color #backgroundColorFormatterNPSgroup {
    thresholds: #7ED251 >=9, #FFBB5C >= 7, #F76373 >= 0,#E0E0E0 <0

  }
  formatter color #backgroundColorFormatterNPS {
    thresholds: #7ED251 >=20, #FFBB5C >= 10, #F76373 <= 10
  }
  formatter color #valueColorFormatter {
    thresholds: #333333 >=9, #333333 >=7, #ffffff >= 0
  }
  formatter color #valueColorFormatterIndex {
    thresholds: #333333 >=8, #333333 >=6, #ffffff >= 0,#E0E0E0 <0
    defaultValue: transparent
  }
  formatter color #valueColorFormatterNPSgroup {
    thresholds: #333333 >=9, #333333 >=7, #ffffff >= 0,#5C5C5C <0
  }
  formatter color #valueColorFormatterNPS {
    thresholds: #333333 >=20, #333333 >=10, #ffffff <= 10
  }
  formatter color #riskTextColorFormatter {
    thresholds: #FFFFFF >= 9, #333333 >= 7,#FFFFFF >=0, #5C5C5C <0
  }
  formatter color #riskTextBgColorFormatter {
    thresholds: #82D854 >= 9,  #F0AD4E >= 7,#FA5263 >=0,#DEDDDD <0
  }
  formatter color #healthTextColorFormatter {
    thresholds: #FFFFFF = 1, #FFFFFF = 2, #333333 = 3,#FFFFFF =4, #333333 =0
  }
  formatter color #healthTextBgColorFormatter {
    thresholds: #82D854 = 1, #D6D854 = 2, #F0AD4E = 3,#FA5263 =4,#cccccc =0
  }
  formatter color #adoptionTextColorFormatter {
    thresholds: #FFFFFF >= 10, #333333 >= 5,#FFFFFF >=0, #333333 < 0
  }
  formatter color #adoptionTextBgColorFormatter {
    thresholds: rgba(126, 210, 81, 0.655) >= 10,  rgba(255, 187, 92, 0.765) >= 5,rgba(247, 99, 114, 0.731) >=0, #cccccc < 0
  }

  //RECODED LABELS
  formatter color #loyaltygroups {
    thresholds: Loyal >= 9, Passive >= 7, Unlikely >= 0
  }
  formatter color #NPSgroups {
    thresholds: Promoter >= 9, Passive >= 7, Detractor >= 0
  }
  formatter color #NPSgroupsContacts {
    thresholds: Silent < 0, Promoter >= 9, Passive >= 7, Detractor >= 0
  }
  formatter color #usertrend {
    thresholds: High >= 10, Med >= 5 , Low >= 0 , Unknown < 0
  }
  formatter color #usagetrend {
    thresholds: Decline < 0, Static >= 5, Growth >=10
  }
  formatter color #adoptionrate {
    thresholds: Low >= 0 , Med >= 5, Active >= 10
  }
  formatter color #spendtrend {
    thresholds: Growth = 10, Static =5, Decline = 0, Unknown <0
  }
  formatter color #LeadScore {
    thresholds: High >= 10, Med >=5, Low >= 0
  }
  formatter color #risklevel {
    thresholds: Low >= 9, Med >=7, High >= 0, Unknown < 0
  }
  formatter color #healthlevel {
    thresholds: Four = 1, One = 4, Two  = 3, Three = 2, Unknown = 0
  }

  //CUSTOM PROPERTIES: FILTER EXPRESSIONS, SEGMENTS, DATE RANGES

  custom properties #filter {

    //CLIENT
    isSent: IIF(respondent:noOfEmailsSent > 0 AND respondent:smtpStatus != "NonDeliveryReport", true, false)
    isResponded: IIF(relationship:status = "complete", true, false)
    isPartial: IIF(relationship:status = "incomplete" AND _IsNull(relationship:Q1) = false, true, false)
    isFailedInvite: IIF((respondent:smtpStatus != "messageSent" AND respondent:smtpStatus != "OptOut") AND respondent:noOfEmailsSent > 0, true, false)
    isNotYetSent: IIF(respondent:noOfEmailsSent = 0, true, false)
    isOptOut: IIF((respondent:OptOut = "3" OR respondent:OptOut = "6") OR respondent:smtpStatus = "OptOut", true, false)
    isClientResponse: IIF(_IsNull(relationship:Q1) = false, true, false)
    isClientSurvey: IIF(clientandteam:combined_sourceid = "p1850259384", true, false)

    //TEAM
    isTeamResponse: IIF(_IsNull(teamcheck:Q1) = false, true, false)
    isTeamSent: IIF(teamcheckresp:noOfEmailsSent > 0 AND teamcheckresp:smtpStatus != "NonDeliveryReport", true, false)
    isTeamSurvey: IIF(clientandteam:combined_sourceid = "p1860215844", true, false)

  }

  //FIXED REPORTING PERIODS
  custom properties #daterange {

//Revenue
    currentPeriodRev: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthRev, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthRev, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthRev, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearRev, true))))
    previousPeriodRev: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.P3MonthRev, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.P6MonthRev, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.P12MonthRev, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.PCalYearRev, true))))


    L3MonthRev: Between(SFDCClosedOpportunities:CloseDate, AddMonth(GetDate(), -3), GetDate()) AND SFDCClosedOpportunities:IsClosed = "true"
    P3MonthRev: Between(SFDCClosedOpportunities:CloseDate, AddMonth(GetDate(), -6), AddMonth(GetDate(), -3)) AND SFDCClosedOpportunities:IsClosed = "true"

    L6MonthRev: Between(SFDCClosedOpportunities:CloseDate, AddMonth(GetDate(), -6), GetDate()) AND SFDCClosedOpportunities:IsClosed = "true"
    P6MonthRev: Between(SFDCClosedOpportunities:CloseDate, AddMonth(GetDate(), -12), AddMonth(GetDate(), -6)) AND SFDCClosedOpportunities:IsClosed = "true"

    L12MonthRev: Between(SFDCClosedOpportunities:CloseDate, AddYear(GetDate(), -1), GetDate()) AND SFDCClosedOpportunities:IsClosed = "true"
    P12MonthRev: Between(SFDCClosedOpportunities:CloseDate, AddYear(GetDate(), -2), AddYear(GetDate(), -1)) AND SFDCClosedOpportunities:IsClosed = "true"


    //to be updated.
    CCalYearRev: InYear(SFDCClosedOpportunities:CloseDate, 0, 0) AND SFDCClosedOpportunities:IsClosed = "true"
    PCalYearRev: InYear(SFDCClosedOpportunities:CloseDate, -1, -1) AND SFDCClosedOpportunities:IsClosed = "true"

    //RELATONSHIP SURVEY
    currentPeriodRel: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthRel, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthRel, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthRel, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearRel, true))))
    previousPeriodRel: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.P3MonthRel, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.P6MonthRel, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.P12MonthRel, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.PCalYearRel, true))))
    currentPeriodRelRate: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthRelRate, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthRelRate, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthRelRate, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearRelRate, true))))
    currentPeriodRelResp: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthRelResp, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthRelResp, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthRelResp, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearRelResp, true))))

    L3MonthRel: Between(relationship:interview_start, AddMonth(GetDate(), -3), GetDate())
    P3MonthRel: Between(relationship:interview_start, AddMonth(GetDate(), -6), AddMonth(GetDate(), -3))
    L3MonthRelRate: Between(relationship:FirstMailedDate, AddMonth(GetDate(), -3), GetDate())
    L3MonthRelResp: Between(respondent:FirstEmailedDate, AddMonth(GetDate(), -3), GetDate())

    L6MonthRel: Between(relationship:interview_start, AddMonth(GetDate(), -6), GetDate())
    P6MonthRel: Between(relationship:interview_start, AddMonth(GetDate(), -12), AddMonth(GetDate(), -6))
    L6MonthRelRate: Between(relationship:FirstMailedDate, AddMonth(GetDate(), -6), GetDate())
    L6MonthRelResp: Between(respondent:FirstEmailedDate, AddMonth(GetDate(), -6), GetDate())

    L12MonthRel: Between(relationship:interview_start, AddYear(GetDate(), -1), GetDate())
    P12MonthRel: Between(relationship:interview_start, AddYear(GetDate(), -2), AddYear(GetDate(), -1))
    L12MonthRelRate: Between(relationship:FirstMailedDate, AddYear(GetDate(), -1), GetDate())
    L12MonthRelResp: Between(respondent:FirstEmailedDate, AddYear(GetDate(), -1), GetDate())

    //to be updated.
    CCalYearRel: InYear(relationship:interview_start, 0, 0)
    PCalYearRel: InYear(relationship:interview_start, -1, -1)
    CCalYearRelRate: InYear(relationship:FirstMailedDate, 0, 0)
    CCalYearRelResp: InYear(respondent:FirstEmailedDate, 0, 0)


    //TEAM CHECK SURVEYM
    currentPeriodTC: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthTC, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthTC, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthTC, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearTC, true))))
    previousPeriodTC: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.P3MonthTC, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.P6MonthTC, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.P12MonthTC, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.PCalYearTC, true))))
    currentPeriodTCRate: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthTCRate, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthTCRate, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthTCRate, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearTCRate, true))))
    currentPeriodTCResp: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthTCResp, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthTCResp, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthTCResp, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearTCResp, true))))

    L3MonthTC: Between(teamcheck:interview_start, AddMonth(GetDate(), -4), GetDate())
    P3MonthTC: Between(teamcheck:interview_start, AddMonth(GetDate(), -7), AddMonth(GetDate(), -4))
    L3MonthTCRate: Between(teamcheck:FirstMailedDate, AddMonth(GetDate(), -4), GetDate())
    L3MonthTCResp: Between(teamcheckresp:FirstEmailedDate, AddMonth(GetDate(), -4), GetDate())

    L6MonthTC: Between(teamcheck:interview_start, AddMonth(GetDate(), -7), GetDate())
    P6MonthTC: Between(teamcheck:interview_start, AddMonth(GetDate(), -13), AddMonth(GetDate(), -7))
    L6MonthTCRate: Between(teamcheck:FirstMailedDate, AddMonth(GetDate(), -7), GetDate())
    L6MonthTCResp: Between(teamcheckresp:FirstEmailedDate, AddMonth(GetDate(), -7), GetDate())

    L12MonthTC: Between(teamcheck:interview_start, AddMonth(AddYear(GetDate(), -1), -1), GetDate())
    P12MonthTC: Between(teamcheck:interview_start, AddMonth(AddYear(GetDate(), -2), -1), AddMonth(AddYear(GetDate(), -1), -1))
    L12MonthTCRate: Between(teamcheck:FirstMailedDate, AddMonth(AddYear(GetDate(), -1), -1), GetDate())
    L12MonthTCResp: Between(teamcheckresp:FirstEmailedDate, AddMonth(AddYear(GetDate(), -1), -1), GetDate())

    CCalYearTC: InYear(teamcheck:interview_start, 0, 0)
    PCalYearTC: InYear(teamcheck:interview_start, -1, -1)
    CCalYearTCRate: InYear(teamcheck:FirstMailedDate, 0, 0)
    CCalYearTCResp: InYear(teamcheckresp:FirstEmailedDate, 0, 0)

    //CASES
    currentPeriodCases: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthCases, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthCases, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthCases, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearCases, true))))
    previousYearCases: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.P3MonthCases, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.P6MonthCases, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.P12MonthCases, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.PCalYearCases, true))))

    L3MonthCases: Between(cases:DateCreated, AddMonth(GetDate(), -3), GetDate())
    P3MonthCases: Between(cases:DateCreated, AddMonth(GetDate(), -6), AddMonth(GetDate(), -3))

    L6MonthCases: Between(cases:DateCreated, AddMonth(GetDate(), -6), GetDate())
    P6MonthCases: Between(cases:DateCreated, AddMonth(GetDate(), -12), AddMonth(GetDate(), -6))

    L12MonthCases: Between(cases:DateCreated, AddYear(GetDate(), -1), GetDate())
    P12MonthCases: Between(cases:DateCreated, AddYear(GetDate(), -2), AddYear(GetDate(), -1))

    CCalYearCases: InYear(cases:DateCreated, 0, 0)
    PCalYearCases: InYear(cases:DateCreated, -1, -1)

   // REL AND TC COMBINED
    currentPeriodTRCom: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthTRCom, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthTRCom, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthTRCom, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearTRCom, true))))
    previousPeriodTRCom: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.P3MonthTRCom, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.P6MonthTRCom, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.P12MonthTRCom, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.PCalYearTRCom, true))))

    L3MonthTRCom: Between(clientandteam:RelationshipSurveyDate, AddMonth(GetDate(), -3), GetDate())
    P3MonthTRCom: Between(clientandteam:RelationshipSurveyDate, AddMonth(GetDate(), -6), AddMonth(GetDate(), -3))

    L6MonthTRCom: Between(clientandteam:RelationshipSurveyDate, AddMonth(GetDate(), -6), GetDate())
    P6MonthTRCom: Between(clientandteam:RelationshipSurveyDate, AddMonth(GetDate(), -12), AddMonth(GetDate(), -6))

    L12MonthTRCom: Between(clientandteam:RelationshipSurveyDate, AddYear(GetDate(), -1), GetDate())
    P12MonthTRCom: Between(clientandteam:RelationshipSurveyDate, AddYear(GetDate(), -2), AddYear(GetDate(), -1))

    CCalYearTRCom: InYear(clientandteam:RelationshipSurveyDate, 0, 0)
    PCalYearTRCom: InYear(clientandteam:RelationshipSurveyDate, -1, -1)

// Finance
    currentPeriodFin: IIF(@timeperiod.selectedOption.label = "Last 3 Months", @daterange.L3MonthFin, IIF(@timeperiod.selectedOption.label = "Last 6 Months", @daterange.L6MonthFin, IIF(@timeperiod.selectedOption.label = "Last 12 Months", @daterange.L12MonthFin, IIF(@timeperiod.selectedOption.label = "Current Calendar Year", @daterange.CCalYearFin, true))))

    L3MonthFin: InQuarter(finance:month, -1, -1)
    L6MonthFin: InQuarter(finance:month, -2, -1)
    L12MonthFin: InQuarter(finance:month, -4, -1)
    CCalYearFin: InYear(finance:month, 0, 0)
  }




  //ELEMENT INDEX SCORES
  custom properties #index {

    NPS: IIF(SFDCAccounts:NPSavg >= 9, 10, IIF(SFDCAccounts:NPSavg >= 7, 5, IIF(SFDCAccounts:NPSavg >= 0, 0)))
    Needs: IIF(SFDCAccounts:NEEDSavg >= 9, 10, IIF(SFDCAccounts:NEEDSavg >= 7, 5, IIF(SFDCAccounts:NEEDSavg >= 0, 0)))
    Value: IIF(SFDCAccounts:VALUEavg >= 9, 10, IIF(SFDCAccounts:VALUEavg >= 7, 5, IIF(SFDCAccounts:VALUEavg >= 0, 0)))
    Relationship: IIF(SFDCAccounts:RELavg >= 9, 10, IIF(SFDCAccounts:RELavg >= 7, 5, IIF(SFDCAccounts:RELavg >= 0, 0)))
    Technology: IIF(SFDCAccounts:TECHavg >= 9, 10, IIF(SFDCAccounts:TECHavg >= 7, 5, IIF(SFDCAccounts:TECHavg >= 0, 0)))

    tNPS: IIF(SFDCAccounts:tNPSavg >= 9, 10, IIF(SFDCAccounts:tNPSavg >= 7, 5, IIF(SFDCAccounts:tNPSavg >= 0, 0)))
    Renew: IIF(SFDCAccounts:RENEWavg >= 9, 10, IIF(SFDCAccounts:RENEWavg >= 7, 5, IIF(SFDCAccounts:RENEWavg >= 0, 0)))
    Benefits: IIF(SFDCAccounts:BENavg >= 9, 10, IIF(SFDCAccounts:BENavg >= 7, 5, IIF(SFDCAccounts:BENavg >= 0, 0)))
    Experience: IIF(SFDCAccounts:EXPavg >= 9, 10, IIF(SFDCAccounts:EXPavg >= 7, 5, IIF(SFDCAccounts:EXPavg >= 0, 0)))

    //CLIENT BEHAVIOUR INDEX SCORES
    SpendTrend: IIF(SFDCAccounts:ltrL12MRev >= 0 OR SFDCAccounts:ltrP12MRev >= 0, IIF(SFDCAccounts:ltrP12MRev = 0, IIF(SFDCAccounts:ltrL12MRev > 0, 5), IIF(SFDCAccounts:revDiff < -10, 0, IIF(SFDCAccounts:revDiff > 10, 10, 5))))
    UserAdoption: IIF(SFDCAccounts:usersLicenses > 0, IIF(SFDCAccounts:usages >= 80, 10, IIF(SFDCAccounts:usages < 40, 0, 5)))
    LeadScore: IIF(count(SFDCMarketLeads:mkto71_Lead_Score) > 0, IIF(average(SFDCMarketLeads:mkto71_Lead_Score) >= 95, 10, IIF(average(SFDCMarketLeads:mkto71_Lead_Score) < 24, 0, 5)))
    ResponseRate: IIF(SFDCAccounts:responseRateL12M >= 50, IIF(SFDCAccounts:noResponsesL12M <= 2, 0, 10), IIF(SFDCAccounts:responseRateL12M >= 0, IIF(SFDCAccounts:noResponsesL12M <= 2, 0, 5)))

  }

  //WEIGHT MODEL
  custom properties #weight {

  //CLIENT FEELING ELEMENTS
    NPS: .05 //Q1
    Needs: .40  //Q12
    Value: .15 //Q3
    Relationship: .10 //Q4
    Technology: .30 //Q7
    //TEAM FEELING ELEMENTS
    tNPS: .05 //Q1
    Renew: .40 //Q2
    Benefits: .15 //Q8
    Experience: .40 //Q9
   //BEHAVIOUR ELEMENTS
    ResponseRate: .10 //Response Rate weight
    LeadScore: .10 //MarketingLeadScore
    SpendTrend: .60 //YoY Revenue
    UserAdoption: .20 //RVA Licensed vs Active
  //FOCUS WEIGHTS
    clientfeeling: .30
    teamfeeling: .30
    doing: .40
  //FOCUS WEIGHTS.SIMPLIFIED
    clientfeeling2: .50
    teamfeeling2: .50

  }

//CALCULATIONS
  custom properties #calculate {
    salesperformance: (Sum(finance:NetsalesquotaachievementAmericasVoC) + Sum(finance:NetsalesquotaachievementAmericasMR) + Sum(finance:NetsalesquotaachievementGlobalVoE) + Sum(finance:NetsalesquotaachievementNordicsVoC) + Sum(finance:NetsalesquotaachievementEMEAVoC) + Sum(finance:NetsalesquotaachievementEMEAMR) + Sum(finance:NetsalesquotaachievementAustralia) + Sum(finance:NetsalesquotaachievementRussia)) / 8 * 100
  }

  //TARGETS
  custom properties #targets {
    // NEED TO CHANGE TO A DYNAMIC
    NPS: 20 // Client NPS
    tNPS: 20 // Internal NPS
    metricAvg: 8
    indexScore: 8
  }

}

//FILTER PANEL
layoutArea toolbar {

  filter hierarchy {
    label: "Sales Organisation"
    hierarchy: hierarchy:21039
    optionLabel: hierarchy:language_text
    smartExpand: true
  }

  filter drillDown {
    drillDown: accountOwner
    label: "Account Owner"
  }

  filter multiselect #AccountTeam {
    label: "Account Team"
    optionsFrom: SFDCAccounts:sAccountTeam
  }

  filter multiselect #clientType {
    label: "Client Type"
    optionsFrom: SFDCAccounts:sClientType
  }

  filter multiselect #industries {
    label: "Industry"
    optionsFrom: SFDCAccounts:Industry
  }

  filter multiselect #typeofcustomer {
    label: "Type of Customer"
    optionsFrom: SFDCAccounts:sTypeOfCustomer
  }
  filter multiselect #riskGroup {
    label: "Risk Priority"
    optionsFrom: SFDCAccounts:riskgroups
  }

  filter multiselect #role {
    label: "Role"
    option checkbox #r1 {
      label: "Decision maker"
      value: contacts:contactRole = "Decision maker"
    }
    option checkbox #r2 {
      label: "Influencer"
      value: contacts:contactRole = "Influencer"
    }
    option checkbox #r3 {
      label: "Champion/Coach"
      value: contacts:contactRole = "Champion/Coach"
    }
    option checkbox #r4 {
      label: "User"
      value: contacts:contactRole = "User"
    }
    option checkbox #r5 {
      label: "Admin/PA"
      value: contacts:contactRole = "Admin/PA"
    }
    option checkbox #r6 {
      label: "Procurement"
      value: contacts:contactRole = "Procurement"
    }
    option checkbox #r7 {
      label: "Other"
      value: contacts:contactRole = "Procurement"
    }
  }

  filter multiselect #annualaccountvalue {
    label: "Revenue - Last 12 Months"
    option checkbox #r1 {
      label: "< $50K"
      value: Between(SFDCAccounts:ltrL12MRev, 1, 50000)
    }
    option checkbox #r2 {
      label: "$50k-$99k"
      value: Between(SFDCAccounts:ltrL12MRev, 50000, 99999.99)
    }
    option checkbox #r3 {
      label: "$100k-$249k"
      value: Between(SFDCAccounts:ltrL12MRev, 100000, 249999.99)
    }
    option checkbox #r4 {
      label: "$250k-$499k"
      value: Between(SFDCAccounts:ltrL12MRev, 250000, 499999.99)
    }
    option checkbox #r5 {
      label: "$500k-$999k"
      value: Between(SFDCAccounts:ltrL12MRev, 500000, 999999.99)
    }
    option checkbox #r6 {
      label: "$1m+"
      value: SFDCAccounts:ltrL12MRev > 999999.99
    }
    option checkbox #r7 {
      label: "No revenue in the last 12 months"
      value: SFDCAccounts:ltrL12MRev <= 0.99 OR _IsNull(SFDCAccounts:ltrL12MRev)
    }

  }


  filter singleselect #timeperiod {
    label: "Time Period"
    canClear: false
    option radio #r1 {
      label: "Last 3 Months"
      value: SFDCAccounts:id != ""
    }
    option radio #r2 {
      label: "Last 6 Months"
      value: SFDCAccounts:id != ""
    }
    option radio #r3 {
      label: "Last 12 Months"
      value: SFDCAccounts:id != ""
      selected: true
    }
    // option radio #r4 {
    //   label: "Current Calendar Year"
    //   value: accounts:id != ""
    // }
  }

  filter singleselect #accountactivitystatus {
    hide: true
    canClear: false
    label: "Account Activity Status"
    option checkbox #r3 {
      label: "Active Client"
      value: SFDCAccounts:accountActivityStatus = "1"
      selected: true
    }
    option checkbox #r4 {
      label: "Inactive Client"
      value: SFDCAccounts:accountActivityStatus = "2"
    }
  }

  filter multiselect #responserate {

    label: "Response Rate - Last 12 Months"
    option checkbox #r1 {
      label: "No Invites sent to contacts"
      value: _IsNull(SFDCAccounts:responseRateL12M)
    }
    option checkbox #r2 {
      label: "Low (<25%)"
      value: SFDCAccounts:responseRateL12M < 25
    }
    option checkbox #r3 {
      label: "OK (>=25%)"
      value: SFDCAccounts:responseRateL12M >= 25
    }
  }


  filter singleselect #voxPopme {
    label: "Voxpopme Filter"

    option checkbox {
      label: "Show Answered Only"
      value: feedback:Q3_vox.answered
    }
    option checkbox {
      label: "Show Skipped Only"
      value: feedback:Q3_vox.skipped
    }
  }

  filter multiselect #storyTheme {
    label: "Story Theme"
    option checkbox {
      label: "Getting you up and running painlessly"
      value: feedback:Q3_vox.answered
    }
    option checkbox {
      label: "Partnership – helping you develop your program over time"
      value: feedback:Q3_vox.answered
    }
    option checkbox {
      label: "Joining up across Customer Journey / Breaking Down Silos / Integration"
      value: feedback:Q3_vox.answered
    }
    option checkbox {
      label: "Business Impact – (Increases in revenue / reduction in costs / driving action)"
      value: feedback:Q3_vox.answered
    }
    option checkbox {
      label: "Driving engagement – Leaders / Front Line"
      value: feedback:q3_vox.answered
    }
    option checkbox {
      label: "Culture Change – becoming more 'customer centric' OR living the client 'Values'"
      value: feedback:Q3_vox.answered
    }
    option checkbox {
      label: "Other"
      value: feedback:Q3_vox.answered
    }
  }
}

page #PortfolioHealth {

  widget search {
    layoutArea: "header"
    source search #ss {
      table: SFDCAccounts:
      value: SFDCAccounts:Name + " (" + SFDCAccounts:Id + ")"
      navigateTo: AccountOverview
    }
  }

  label: "Account Health"
  widget summary {
    size: large

    infobox {
      label: "Top Level Summary"
      info: "Overall Assessment of risk of portfolio defined by the applied hierarchy filter. Calculated as a weighted index as illustrated by Risk Modeller graphic below., incorporating

 - **Client Feeling:**  Currently measured by Relationship Survey NPS only

- **Client Behaviour:** Currently measured by Spend Trend, Product Usage, Response Rate, Marketing Engagement

- **Team Feeling:** Currently measured by Account Manager perception of NPS"
    }

    tile risk {
      label: "Portfolio Risk Priority"
      showThermometer: false

      value: average(SFDCAccounts:overallIndex)
      textValue: IIF(_IsNull(average(SFDCAccounts:overallIndex)), "Unknown", IIF(average(SFDCAccounts:overallIndex) >= 8, "Priority 4", IIF(average(SFDCAccounts:overallIndex) >= 6, "Priority 3", "Priority 2")))

      min: 0
      max: 5

      target: @targets.indexScore

   //   renewal: first(SFDCAccounts:AccountRenewalDate, SFDCAccounts:AccountRenewalDate, InMonth(SFDCAccounts:AccountRenewalDate, 1, 36))
      revenue: sum(SFDCAccounts:ltrL12MRev)
      revenueLabel: "Last 12 mnths Rev"
    }
    tile metric {
      label: "Client Behaviour"
      value: round(average(SFDCAccounts:clientBehaviourIndex), 1)
      target: @targets.indexScore
    }
    tile metric {
      label: "Client Feeling"
      value: round(average(SFDCAccounts:clientFeelingIndex), 1)
      target: @targets.indexScore

    }
    tile metric {
      label: "Team Feeling"
      value: round(average(SFDCAccounts:teamFeelingIndex), 1)
      target: @targets.indexScore
    }
  }
  widget markdown {

    infobox {
      label: "Decision Modeller"
      info: "**Client Feeling**

**Currently measured by Relationship Survey only**
- NPS (5%)
- Fulfils my Needs (40%)
- Delivers value to my organisation (15%)
- Satisfaction with the team (10%)
- Satisfaction with the technology (30%)
 *We will incorporate Implementation, Support & Training surveys into this metric*

**Client Behavior**

- Spend Trend = Change in revenue in last 12 months
- Product Usage = RVA's used compared to those sold
- Response Rate = For Relationship survey only,
- Marketing Engagement = Index based on data available in SFDC
    - **Usage does not include usage of RVAs for Active Dashboards**

**Team Feeling**

*Currently measured by Account Manager perception of *

- NPS (5%)
- Liklihood to renew (40%)
- Recognise benefits across the organisation (15%)
- Confirmit support experience (40%)
"
    }

    size: small
    label: "Decision Modeller"
    markdown: "
![Risk Factors](http://survey.euro.confirmit.com/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/EMPOWER/Risk%20Modeller.PNG)
"
  }

  //WIDGET NOT WORKING - CANNOT HAVE MULTIPLE SOURCES ON ONE CHART WHERE SOME SOURCES DO NOT HAVE DIRECT
  //RELATIONSHIPS WITH EACH OTHER.
  widget chart {

    infobox {
      label: "Risk Trend"
      info: "**NOTE:** Currently we can only show Client Feeling score due to limitation in Studio.

- We will add other trend lines as soon as soon as available"
    }

    filter expression {
      value: @daterange.currentPeriodRel
    }

    label: "Risk Trend"
    //  //palette: "#2B3E50","#DF691A","#4bf442"
    // palette: "#2B3E50","#54bc23"
    size: medium
    legend: bottomCenter
    gridLines: none
    removeEmptyCategories: true

    // chart area {
    //   lineType: monotone
    // }

    chart line {
      //lineType: basis
      dotSize: 5

    }

    series #ss1 {
      value: round(average(SFDCAccounts:clientBehaviourIndex), 1)
     // format: onedecimal
      label: "Client Behaviour"
    }
    series #ss2 {
      value: round(average(SFDCAccounts:clientFeelingIndex), 1)
    //  format: onedecimal
      label: "Client Feeling"

    }
    series #ss3 {
      value: round(average(SFDCAccounts:teamFeelingIndex), 1)
   //   format: onedecimal
      label: "Team Feeling"
    }

    series #ss4 {
      value: round(average(SFDCAccounts:overallIndex), 1)
      //format: onedecimal
      label: "Overall"
      chart line {
        lineType: linear
        dotSize: 0
        lineWidth: 5
      }
    }

    category overlappingDate {
      value: relationship:interview_start
      breakdownBy: calendarMonth
      start: "-13 months"
      end: "0 days"
      startShift: "-12 months"
      endShift: "0 months"
      format: monthlabel
    }
  }
  widget responseRate {

    infobox {
      label: "Feedback Response Rate"
      info: "The Feedback Response Rate widget provides a breakdown of the possible response categories for the relationship survey for the time period selected (default last 12 month rolling).
      *Click on a bar to provide a list of clients*"
    }

    size: small
    label: "Feedback Response Rate"

    table: respondent:
    rem
    tile statuses {
      breakBy: respondent:responseStatus
      value: count(respondent:responseStatus, @daterange.currentPeriodRelResp)
      chart: "bar"
      palette: '#CCCCCC', '#f44245', '#f49541','#f4ee41','#82D854'
      //format:
      percentFormat: percentage
      navigateTo: "Response Management"
    }

    //ISSUE HERE - WHY IS IT NOT TAKING THE RIGHT COUNTS FOR NO EMAILED
    tile value {
      label: "Invitations Delivered"
      value: count(respondent:respid, @daterange.currentPeriodRelResp AND @filter.isSent)
      //format: responsesFormat
    }
    tile value {
      label: "Response rate"
      format: percentage
      value: count(relationship:responseid, (@filter.isResponded OR @filter.isPartial) AND @daterange.currentPeriodRelRate) * 100 / count(respondent:respid, @daterange.currentPeriodRelResp AND @filter.isSent) // invite sent in 2018
    }
  }




  widget chart #revenuerisk {


    filter expression {
      value: InMonth(SFDCAccounts:AccountRenewalDate, 0, 6)
    }
    infobox {
      label: "Revenue Risk 6mth Forecast"
      info: "Breakdown of portfolio by month and risk level.
      **Value:** Sum of closed opportunities for the last 12 months"
    }

    palette: #FA5263,#F0AD4C,#D6D854,#82D854,#cccccc
    table: SFDCAccounts:

    label: "Revenue Risk - 6mth Forecast"
    size: medium
    navigateTo: "Accounts in Segment"
    legend: bottomCenter

    chart bar {
      dataLabel: valueThenPercent
      mode: stacked
    }
    series {
      value: sum(SFDCAccounts:ltrL12MRev)
      format: UScurrency
      breakdownBy cut {
        value: SFDCAccounts:riskgroups
      }
    }
    category date {
      value: SFDCAccounts:AccountRenewalDate
      breakdownBy: calendarMonth
      format: monthlabel
      start: "0 months"
      end: "6 months"
      removeEmpty: true
    }
    removeEmptyCategories: true
    axis primary {
      format: UScurrency
    }

    base {
      value: count(SFDCAccounts:riskgroups)
    }

  }



  widget chart #barAlertTypeByStatus {

    infobox {
      label: "Alert Type by Status"
      info: "Overview of type of alerts by status. Click on a category to provide a list of cases."
    }
    table: cases:
    legend: bottomCenter

    filter expression {
      value: @daterange.currentPeriodCases
      filtertype: "preAggregate"
    }
    //palette: #F51010,#EEAE25,#FFED48,#B22E02,#1EC210,#CCCCCC,#000000
    label: "Alert Type by Status"
    size: medium

    format: nodecimal
    navigateTo: "Customer Alerts"

    chart bar {
      stacked: true
    }
    series {
      value: count(cases:Workflow)
      breakdownBy cut {
        value: cases:lk_1545
      }
    }
    category cut {
      value: cases:Workflow
    }
    base {
      value: count(cases:Workflow)
    }
  }

  widget accountList {

    infobox {
      label: "Account Risk"
      info: "Full breakdown of the KPIs for all Active Clients with drill down available to individual Accounts

**Lifetime Value:** All closed opportunities

**Spend Trend:** Change in Revenue Last 12 mths compared to Previous 12 mths

**Overall Risk:** Index combinging Client & Team Feeling and Client Behavior

**Behavior Risk:**

- Spend Trend = Change in revenue in last 12 months
- Product Usage = RVA's used compared to those sold
- Response Rate = For Relationship survey only ,
- Marketing Engagement = Index based on data available in SFDC

**Client Feeling Risk:**

- Avg Relationship Survey NPS for the last 12 months

**Team Feeling Risk:**

- Latest NPS score from the Account Healthcheck completed by Account Manager

**Last Invites and Response:** Client Relationship survey only at this time

**Last Team Check:** Completed by Account Manager"
    }

    label: "Account Risk"
    table: SFDCAccounts:
    sortColumn: noresponsel12M
    sortOrder: descending
    navigateTo: AccountOverviewModal
    size: large
    take: 50
    paginationType: paging
    rowsPerPage: 50,100,150
    headerNumberOfLines: 4


    view metric #risklevel {
      backgroundColorFormatter: riskTextBgColorFormatter
      valueColorFormatter: riskTextColorFormatter
      Size: small
    }

    view metric #healthlevel {
      backgroundColorFormatter: healthTextBgColorFormatter
      valueColorFormatter: healthTextColorFormatter
      Size: small
    }

    view metric #riskformat {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    view metric #adoptionlevelbehaviour {
      backgroundColorFormatter: adoptionTextBgColorFormatter
      valueColorFormatter: adoptionTextColorFormatter
      fontSize: small
    }
    // column link {
    //   label: "Horizons Info"
    //   value: "view"
    //   link href {
    //     address: "https://studio.euro.confirmit.com/apps/dashboard/2898/accountHorizonsInfo?expr=fromcrmconnector.SFDCAccounts_v6_0_1&selected=" + ToText(SFDCAccounts:id)
    //   }

    // }
    column value #account {
      label: "Account"
      value: SFDCAccounts:Name
      rowHeader: true
      enableColumnFilter: true
    }

    column value #noresponsel12M {
      label: "# Responses L12M"
      value: SFDCAccounts:noresponsesL12M
      format: nodecimal
      align: right
    }
    column metric #risk {
      label: "Overall Risk Priority"
      value: IIF((SFDCAccounts:clientFeelingRiskCategory = "High" AND SFDCAccounts:clientBehaviourRiskCategory = "High") AND (SFDCAccounts:teamFeelingRiskCategory = "High" OR SFDCAccounts:teamFeelingRiskCategory = "Unknown"), 4, IIF(_IsNull(SFDCAccounts:overallIndex), 0, IIF(SFDCAccounts:overallIndex >= 8, 1, IIF(SFDCAccounts:overallIndex >= 6, 2, 3))))
      align: center
      format: healthlevel
      view: healthlevel
      target: 10
    }
    column metric #behaviourlabel {
      label: "Behaviour Risk"
      value: IIF(SFDCAccounts:clientBehaviourIndex >= 0, SFDCAccounts:clientBehaviourIndex, -1)
      align: center
      format: risklevel
      view: risklevel
      target: 8
    }
    column metric #spendtrend {
      label: "Spend Trend"
      value: IIF(@index.SpendTrend >= 0, @index.SpendTrend, -1)
      format: spendtrend
      target: 10
      align: center
      view: adoptionlevelbehaviour
    }
    column value #revL12M {
      label: "Last 12 mths Rev"
      value: SFDCAccounts:ltrL12MRev
      format: UScurrency
      align: right
    }
    column value #revP12M {
      label: "Prev 12 mths Rev"
      value: SFDCAccounts:ltrP12MRev
      format: UScurrency
      align: right
    }

    column value #totalAccountValue {
      label: "Lifetime Value"
      value: SFDCAccounts:TotalAccountValue_USD
      format: UScurrency
      align: right
    }

    column metric #cfeeling2label {
      label: "Client Feeling Risk"
      value: IIF(SFDCAccounts:clientFeelingIndex >= 0, SFDCAccounts:clientFeelingIndex, -1)
      align: center
      format: risklevel
      view: risklevel
      target: 8
    }
    column value #noInvitesL12M {
      label: "# Invites L12M"
      value: SFDCAccounts:invitedL12M
      align: center
    }
    column value #LastInvite {
      label: "Last Invite Sent"
      value: last(respondent:smtpStatusDate, respondent:smtpStatusDate, @filter.isSent)
      format: dateDefaultFormatter
      align: center
    }
    column value #LastResponse {
      label: "Last Response"
      value: last(relationship:interview_start, relationship:interview_start, @filter.isPartial OR @filter.isResponded)
      format: dateDefaultFormatter
      align: center
    }
    column metric #tfeeling2label {
      label: "Team Feeling Risk"
      value: iif(SFDCAccounts:teamFeelingIndex >= 0, SFDCAccounts:teamFeelingIndex, -1)
      align: center
      format: risklevel
      view: risklevel
      target: 10
    }
    column value #LastTeamCheckInvite {
      label: "Last Team Check Sent"
      value: last(teamcheckresp:smtpStatusDate, teamcheckresp:smtpStatusDate, @filter.isTeamSent)
      format: dateDefaultFormatter
      align: center
    }
    column value #LastTeamCheckResponse {
      label: "Last Team Check Response"
      value: last(teamcheck:interview_start, teamcheck:interview_start, _IsNull(teamcheck:Q1) = false)
      format: dateDefaultFormatter
      align: center
    }
  }
}

page #AccountsinSegment {

  modal: true
  label: "Accounts in segment"

  widget title {
    tile value {
      value: @pageFilters.summaryText
    }
  }

  widget accountList {

    infobox {
      label: "Account Risk"
      info: "The Account Risk widget provides a list of accounts that fit within the filtered portfolio along with their risk calculation and scores associated with the dimensions that comprise this score. The risk calculation is a weighted index that examines the customers feelings as measured by our Empower program, behavior measured through our financial and Salesforce data, and our alignment with their feelings as measured by our VoCe program. Clicking on an account will open the Account Overview page for that specific account."
    }

    label: "Account Risk"
    table: SFDCAccounts:
    sortColumn: account
    sortOrder: ascending
    navigateTo: AccountOverviewModal
    size: large

    view metric #risklevel {
      backgroundColorFormatter: riskTextBgColorFormatter
      valueColorFormatter: riskTextColorFormatter
      Size: small
    }

    view metric #healthlevel {
      backgroundColorFormatter: healthTextBgColorFormatter
      valueColorFormatter: healthTextColorFormatter
      Size: small
    }

    view metric #riskformat {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    view metric #adoptionlevelbehaviour {
      backgroundColorFormatter: adoptionTextBgColorFormatter
      valueColorFormatter: adoptionTextColorFormatter
      fontSize: small
    }
    column value #account {
      label: "Account"
      value: SFDCAccounts:Name
      rowHeader: true
    }
    column metric #risk {
      label: "Overall Risk"
      value: IIF((SFDCAccounts:clientFeelingRiskCategory = "High" AND SFDCAccounts:clientBehaviourRiskCategory = "High") AND (SFDCAccounts:teamFeelingRiskCategory = "High" OR SFDCAccounts:teamFeelingRiskCategory = "Unknown"), 4, IIF(_IsNull(SFDCAccounts:overallIndex), 0, IIF(SFDCAccounts:overallIndex >= 8, 1, IIF(SFDCAccounts:overallIndex >= 6, 2, 3))))
      align: center
      format: healthlevel
      view: healthlevel
      target: 10
    }
    column metric #behaviourlabel {
      label: "Behaviour Risk"
      value: IIF(SFDCAccounts:clientBehaviourIndex >= 0, SFDCAccounts:clientBehaviourIndex, -1)
      align: center
      format: risklevel
      view: risklevel
      target: 8
    }
    column metric #spendtrend {
      label: "Spend Trend"
      value: IIF(@index.SpendTrend >= 0, @index.SpendTrend, -1)
      format: spendtrend
      target: 10
      align: center
      view: adoptionlevelbehaviour
    }
    column value #revL12M {
      label: "Last 12 mths Rev"
      value: SFDCAccounts:ltrL12MRev
      format: UScurrency
      align: right
    }
    column value #revP12M {
      label: "Prev 12 mths Rev"
      value: SFDCAccounts:ltrP12MRev
      format: UScurrency
      align: right
    }

    column value #totalAccountValue {
      label: "Lifetime Value"
      value: SFDCAccounts:TotalAccountValue_USD
      format: UScurrency
      align: right
    }

    column metric #cfeeling2label {
      label: "Client Feeling Risk"
      value: IIF(SFDCAccounts:clientFeelingIndex >= 0, SFDCAccounts:clientFeelingIndex, -1)
      align: center
      format: risklevel
      view: risklevel
      target: 8
    }
    column value #noInvitesL12M {
      label: "# Invites L12M"
      value: SFDCAccounts:invitedL12M
      align: center
    }
    column value #LastInvite {
      label: "Last Invite Sent"
      value: last(respondent:smtpStatusDate, respondent:smtpStatusDate, @filter.isSent)
      format: dateDefaultFormatter
      align: center
    }
    column value #LastResponse {
      label: "Last Response"
      value: last(relationship:interview_start, relationship:interview_start, @filter.isPartial OR @filter.isResponded)
      format: dateDefaultFormatter
      align: center
    }
    column metric #tfeeling2label {
      label: "Team Feeling Risk"
      value: iif(SFDCAccounts:teamFeelingIndex >= 0, SFDCAccounts:teamFeelingIndex, -1)
      align: center
      format: risklevel
      view: risklevel
      target: 10
    }
    column value #LastTeamCheckInvite {
      label: "Last Team Check Sent"
      value: last(teamcheckresp:smtpStatusDate, teamcheckresp:smtpStatusDate, @filter.isTeamSent)
      format: dateDefaultFormatter
      align: center
    }
    column value #LastTeamCheckResponse {
      label: "Last Team Check Response"
      value: last(teamcheck:interview_start, teamcheck:interview_start, _IsNull(teamcheck:Q1) = false)
      format: dateDefaultFormatter
      align: center
    }
  }
}

page account #AccountOverviewModal {
  label: "Account Overview"

  modal: true

  mainTable: SFDCAccounts:

  widget title {
    table: SFDCAccounts:

    layout column {
      layout row {
        layout column {
          tile value #c {
            value: SFDCAccounts:Name
          }

        }
        layout column {
          tile role {
            value: SFDCAccounts:AccountOwnerName
          }
        }
        layout column {
          tile company {
            value: SFDCAccounts:SalesRegion
          }
        }
      }
      layout row {
        tile company {
          value: "ID: " + ToText(SFDCAccounts:id)
        }
      }
      layout row {
        tile company {
          value: "Earliest Renewal Date: " + Left(ToText(SFDCAccounts:AccountRenewalDate), 10)
        }
      }
      layout row {
        tile company {
          value: "Renewals: " + SFDCAccounts:Agreement_Last_Dates
        }
      }
      // layout row {
      //   tile company {
      //     value: "On-Premise Renewal: " + ToText(CalendarDate(SFDCAccounts:AccountRenewalDateOnPremise))
      //   }
      //}
    }
  }
  widget summary {

    infobox {
      label: "Overall Risk Summary"
      info: "The top level summary widget provides a quick view of the current performance within the dimensions used to identify level of risk for the selected account. The Risk calculation is a weighted index that examines the customer's feelings (as measured by our Empower program), behavior (measured through our financial and Salesforce data), and our alignment with their feelings (as measured by our VoCe program)."
    }

    size: large
    table: SFDCAccounts:

    tile risk {
      label: "Overall Risk"
      showThermometer: false
      value: SFDCAccounts:overallIndex
      textValue: SFDCAccounts:overallHealthRiskCategory
      min: 0
      max: 10
      target: @targets.indexScore
      //renewal: SFDCAccounts:AccountRenewalDate
      revenue: SFDCAccounts:ltrL12MRev
      revenueLabel: "Last 12 mnths Rev"

    }
    tile metric {
      label: "Client Behaviour"
      value: SFDCAccounts:clientBehaviourIndex
      target: @targets.indexScore
    }
    tile metric {
      label: "Client Feeling"
      value: SFDCAccounts:clientFeelingIndex
      target: @targets.indexScore
    }

    tile metric {
      label: "Team Feeling"
      value: SFDCAccounts:teamFeelingIndex
      target: @targets.indexScore
    }
    tile casesStatus {
      open: count(cases:CaseId)
      overdue: count(cases:overdue, cases:overdue = "Yes")
    }
    tile casesStatus {
      label: "Open Support tickets"
      open: sum(TicketSummary:count, TicketSummary:StatusId = 1)
      overdue: sum(TicketSummary:count, TicketSummary:StatusId = 1)
      showOverdueText: false

    }
  }

  widget contactList {
    label: "Account Contacts: Latest Response"
    infobox {
      label: "Account Contacts: Latest Response"
      info: "The Contacts widget provides a list of all contacts currently associated with this account within Salesforce."
    }

    view metric #npsgroup {
      backgroundColorFormatter: backgroundColorFormatterNPSgroup
      valueColorFormatter: valueColorFormatterNPSgroup
    }

    table: contacts:
    sortColumn: lastResponse
    sortOrder: descending
    size: large
    navigateTo: "Contact Overview"

    column value #name {
      label: "Name"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }
    // column value #country {
    //   label: "Country"
    //   value: contacts:MailingCountry
    // }
    column date #lastResponse {
      label: "Last Feedback Date"
      value: last(relationship:interview_start, relationship:interview_start, _IsNull(relationship:Q1) = false)
      align: center
    }
    column metric #nps {
      label: "NPS Group"
      value: IIF(last(score(relationship:Q1), relationship:interview_start, _IsNull(relationship:Q1) = false) >= 0, last(score(relationship:Q1), relationship:interview_start, _IsNull(relationship:Q1) = false), -1)
      align: center
      view: npsgroup
      target: 9
      format: NPSgroupsContacts
    }
    column date #lastInvited {
      label: "Last Invite Date"
      value: last(respondent:smtpStatusDate, respondent:smtpStatusDate)
      align: center
    }
    column value #comments {
      label: "Recent Comment"
      value: last(relationship:Q2, relationship:interview_start, _IsNull(relationship:Q1) = false)
    }

    column value #noCases {
      label: "Total Cases"
      value: count(cases:CaseId)
      align: center
    }

    column value #overdueCases {
      label: "Overdue Cases"
      value: count(cases:CaseId, cases:overdue = "Yes")
      align: center
    }

  }

  widget dataGridBeta #clientBehaviourSummary {
    label: "Client Behaviour (Last 12 months)"
    size: small

    // suppressRule {
    //   criteria: COUNT(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRel) = 0
    //   label: "No responses to the relationship survey in the last 12 months"
    // }

    infobox {
      label: "Client Behaviour"
      info: "The Client Behaviour widget provides a view of all of the operational level data used to determine the overall Client Behavior score.

**Client Behavior**

- Spend Trend = Change in revenue in last 12 months
- Product Usage = RVA's used compared to those sold
- Response Rate = For Relationship survey only,
- Marketing Engagement = Index based on data available in SFDC
    - **Usage does not include usage of RVAs for Active Dashboards**"
    }

    view comparativeStatistic #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
    }

    view comparativeStatistic #adoptionlevelbehaviour {
      backgroundColorFormatter: adoptionTextBgColorFormatter
      valueColorFormatter: adoptionTextColorFormatter
    }

    view comparativeStatistic #index {
      backgroundColorFormatter: backgroundColorFormatterIndex
      valueColorFormatter: valueColorFormatterIndex
    }

    row {
      //label: "Client Feeling"

    }
    column {
      label: "Client Behav."
      cell {
        value: iif(SFDCAccounts:clientBehaviourIndex >= 0, SFDCAccounts:clientBehaviourIndex, -1)
        target: 8
        view: index
      }
    }
    column {
      label: "User Adopt."
      cell {
        value: IIF(@index.UserAdoption >= 0, @index.UserAdoption, -1)
        format: usertrend
        view: adoptionlevelbehaviour
        target: 10
      }
    }
    column {
      label: "RVA used / purch."
      cell {
        value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)"))
      }
    }
    column {
      label: "Mrkt Eng."
      cell {
        value: @index.LeadScore
        format: LeadScore
        view: adoptionlevelbehaviour
        target: 10
      }

    }
    column {
      label: "# Mrkt Contacts"
      cell {
        value: count(SFDCMarketLeads:Id)
        format: nodecimal
        align: center
      }
    }
    column {
      label: "Response Rate"
      cell {
        value: SFDCAccounts:responseRateL12M
        format: percentage
        align: center
      }
    }
    column {
      label: "Spend Trend"
      cell {
        value: @index.SpendTrend
        format: spendtrend
        view: adoptionlevelbehaviour
        target: 10
      }
    }
    column {
      label: "Rev. Diff (%)"
      cell {
        value: SFDCAccounts:revDiff
        //format: percentageonedecimal
        align: right
      }
    }
    column {
      label: "Last 12Mth Rev."
      cell {
        value: SFDCAccounts:ltrL12MRev
        format: UScurrency
        align: right
      }
    }
    column {
      label: "Prev 12Mth Rev."
      cell {
        value: SFDCAccounts:ltrP12MRev
        format: UScurrency
        align: right
      }
    }
    column {
      label: "Future - Best Case / Closed / Commit / Pipeline"
      cell {
        value: SFDCAccounts:FutureBCCCP
        format: UScurrency
        align: right
      }
    }

  }

  widget dataGridBeta #clientFeelingSummary {
    label: "Client feeling (Last 12 months average)"
    size: small

    // suppressRule {
    //   criteria: COUNT(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRel) = 0
    //   label: "No responses to the relationship survey in the last 12 months"
    // }

    infobox {
      label: "Client Feeling"
      info: "The Client Feeling widget provides a consolidated view of the survey questions/responses from the Client Relationship and Implementation surveys that are currently being used to determine the Client Feeling score.

**Currently measured by Relationship Survey only**
- NPS (5%)
- Fulfils my Needs (40%)
- Delivers value to my organisation (15%)
- Satisfaction with the team (10%)
- Satisfaction with the technology (30%)
 *We will incorporate Implementation, Support & Training surveys into this metric*"
    }

    view comparativeStatistic #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
    }

    view comparativeStatistic #index {
      backgroundColorFormatter: backgroundColorFormatterIndex
      valueColorFormatter: valueColorFormatterIndex
      fontsize: large
    }

    row {
      //label: "Client Feeling"
    }

    column {
      label: "Client Feeling"
      cell {
        value: iif(SFDCAccounts:clientFeelingIndex >= 0, SFDCAccounts:clientFeelingIndex, -1)
        target: 8
        view: index
      }
    }
    column {
      label: "# Responses"
      cell {
        value: COUNT(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRel)
        format: integerDefaultFormatter
      }
    }
    column {
      label: "Likelihood to recommend"
      cell {
        value: iif(SFDCAccounts:NPSavg >= 0, SFDCAccounts:NPSavg, -1)
        target: 9
        view: metric
      }

    }
    column {
      label: "Support Business Needs"
      cell {
        value: iif(SFDCAccounts:NEEDSavg >= 0, SFDCAccounts:NEEDSavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Added Value"
      cell {
        value: iif(SFDCAccounts:VALUEavg >= 0, SFDCAccounts:VALUEavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Relationship Satisfaction"
      cell {
        value: iif(SFDCAccounts:RELavg >= 0, SFDCAccounts:RELavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Technology Satisfaction"
      cell {
        value: iif(SFDCAccounts:TECHavg >= 0, SFDCAccounts:TECHavg, -1)
        target: 9
        view: metric
      }
    }
  }

  widget dataGridBeta #teamFeelingSummary {

    // suppressRule {
    //   criteria: count(teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC) = 0
    //   label: "No responses to the team check survey in the last 12 months"
    // }

    infobox {
      label: "Team Feeling"
      info: "The Team Feeling widget provides a consolidated view of the survey questions/responses from the latest internal Health Check (and Implementation surveys - TBC) used to determine the Team Feeling score.

**Team Feeling**

*Currently measured by Account Manager perception of *

- NPS (5%)
- Liklihood to renew (40%)
- Recognise benefits across the organisation (15%)
- Confirmit support experience (40%)"
    }

    label: "Team feeling (Latest response in last 12 months)"
    size: small

    view comparativeStatistic #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small

    }
    view comparativeStatistic #index {
      backgroundColorFormatter: backgroundColorFormatterIndex
      valueColorFormatter: valueColorFormatterIndex
    }
    row {
      //label: "Client Feeling"

    }
    column {
      label: "Team Feeling"
      cell {
        value: iif(SFDCAccounts:teamFeelingIndex >= 0, SFDCAccounts:teamFeelingIndex, -1)
        target: 8
        view: index
      }
    }
    column {
      label: "Latest Response Received (L12 Months)"
      cell {
        value: last(teamcheck:interview_start, teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC)
        format: dateDefaultFormatter

      }
    }
    column {
      label: "Likelihood to recommend"
      cell {
        value: iif(SFDCAccounts:tNPSavg >= 0, SFDCAccounts:tNPSavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Likelihood To Renew"
      cell {
        value: iif(SFDCAccounts:RENEWavg >= 0, SFDCAccounts:RENEWavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Recognises benefits"
      cell {
        value: iif(SFDCAccounts:BENavg >= 0, SFDCAccounts:BENavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Confirmit support experience"
      cell {
        value: iif(SFDCAccounts:EXPavg >= 0, SFDCAccounts:EXPavg, -1)
        target: 9
        view: metric
      }
    }

  }


  widget contactList {

    infobox {
      label: "Team Checks"
      info: "TBC."
    }

    label: "Team Check: History"

    table: teamcheck:
    sortColumn: lastResponse
    sortOrder: descending
    size: large

    navigateTo: TeamCheckResponse


    view metric #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
    }

    view metric #npsgroup {
      backgroundColorFormatter: backgroundColorFormatterNPSgroup
      valueColorFormatter: valueColorFormatterNPSgroup
    }

    column value #name {
      label: "Name"
      value: teamcheck:AccountOwner
    }

    column date #lastInvited {
      label: "Invite Date"
      value: teamcheck:FirstMailedDate
      align: center
    }

    column date #lastResponse {
      label: "Feedback Date"
      value: teamcheck:interview_start
      align: center
    }
    column metric #nps {
      label: "NPS Group"
      value: score(teamcheck:Q1)
      view: npsgroup
      target: 9
      align: center
      format: NPSgroupsContacts
    }

    column metric #ltr {
      label: "Recommend"
      value: score(teamcheck:Q1)
      align: center
      target: 9
      view: metric
    }

    column metric #renew {
      label: "Renew"
      value: score(teamcheck:Q2)
      align: center
      target: 9
      view: metric
    }

    column metric #recognise {
      label: "Benefits"
      value: score(teamcheck:Q8)
      align: center
      target: 9
      view: metric
    }

    column metric #supportexerience {
      label: "Support"
      value: score(teamcheck:Q9)
      align: center
      target: 9
      view: metric
    }
  }

  widget dataGridBeta #Opportunities2 {
    label: "Last 24 Months Rolling & Future Opportunities"
    size: large

    filter expression {
      value: (Between(SFDCClosedOpportunities:CloseDate, AddYear(GetDate(), -2), GetDate()) AND SFDCClosedOpportunities:IsClosed = "true") OR SFDCClosedOpportunities:CloseDate > GetDate()
    }

    row cut {
      value: SFDCClosedOpportunities:Name + " (" + SFDCClosedOpportunities:Id + ")"
      total: none

    }

    column {
      label: "Opportunity Closed Date"

      cell {

        value: Max(SFDCClosedOpportunities:CloseDate)
        format: dateDefaultFormatter
      }
    }
    column {
      label: "Opportunity Status"

      cell {
        value: Max(SFDCClosedOpportunities:ForecastCategoryName)
      }
    }
    column {
      label: "Opportunity Amount ($)"
      cell {
        value: Sum(SFDCClosedOpportunities:Amount_USD)
        format: UScurrency
      }
    }
  }


  widget chart #eJournalTicketCategories {
    label: "Support Tickets by Category (last 12 months)"
    size: medium
    legend: topCenter
    layout: vertical

    chart bar {
      mode: stacked
      dataLabel: valueThenPercent
    }
    series {
      value: sum(TicketSummary:count)
      breakdownBy cut {
        value: IIF(TicketSummary:StatusId = 2, "Closed Tickets", "Open Tickets")
      }
    }
    category cut #categoryName {
      value: TicketCategories:fullname
      label: "Ticket Categories"
    }
    axis category {
     // orientation: 90
    }

    margin {
      //bottom: 120
      left: 200
    }
    axis primary {
      //axisLine: false

    }
  }

  widget markdown {
    label: " "
    markdown: "- Please note that the initial mapping of SFDC Acounts to Horizons accounts were done manually so there may be a small % of accounts that are unmapped or mapped incorrectly.
    - Only On-Demand usage data is currently included.
    - Additionally the usage data e.g. number RVAs used vs purchased, is not complete because usage data is not available for all products in Horizons, only Reportal and Dashboard / Instant Analytics is covered in the results."

    size: large

  }

  widget contactSurveyResponse {
    label: "Horizons Information"
    size: large
    table: SFDCAccounts:

    tab {
      label: "SITES SUMMARY"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Sites"
          value: ToText("EURO:" + IIF(count(usageAccounts:Id, usageAccounts:site = "euro") > 0, "YES", "No") + " / US:" + IIF(count(usageAccounts:Id, usageAccounts:site = "us") > 0, "YES", "No") + " / AUS:" + IIF(count(usageAccounts:Id, usageAccounts:site = "aus") > 0, "YES", "No") + " /CA:" + IIF(count(usageAccounts:Id, usageAccounts:site = "ca") > 0, "YES", "No") + " / HK:" + IIF(count(usageAccounts:Id, usageAccounts:site = "hk") > 0, "YES", "No"))
        }
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id)
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize)
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize)
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData)
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData)
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData)
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate())
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate())
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52) > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51) > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56) > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3) > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55) > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20) > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37) > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49) > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63) > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34) > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61) > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57) > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39) > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44) > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25) > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62) > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54) > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28) > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53) > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21) > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7) > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29) > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64) > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8) > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27) > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33) > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16) > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40) > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48) > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24) > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2) > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46) > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60) > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59) > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58) > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45) > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50) > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22) > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22) > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives") > 0, "YES", "No")
        }

      }

    }

    tab {
      label: "EUROPE"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "euro")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "euro")
          format: nodecimal
        }

        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "euro")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "euro")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "euro")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "euro")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "USA"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "us")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "us")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "us")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "us")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "us")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "AUSTRALIA"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "aus")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "aus")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "aus")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "aus")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "aus")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "CANADA"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "ca")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "ca")
          format: nodecimal
        }

        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "ca")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "ca")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "ca")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "ca")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "HONG KONG"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "hk")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "hk")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "hk")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "hk")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "hk"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "hk")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "hk")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "hk"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "hk")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "hk")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
      }
    }

  }
}

page account #AccountOverview {
  label: "Account Overview"

  hide: true

  widget search {
    layoutArea: "header"
    source search #ss2 {
      table: SFDCAccounts:
      value: SFDCAccounts:Name + " (" + SFDCAccounts:Id + ")"
      navigateTo: AccountOverview
    }
  }

  mainTable: SFDCAccounts:

  widget title {
    table: SFDCAccounts:

    layout column {
      layout row {
        layout column {
          tile value #c {
            value: SFDCAccounts:Name
          }

        }
        layout column {
          tile role {
            value: SFDCAccounts:AccountOwnerName
          }
        }
        layout column {
          tile company {
            value: SFDCAccounts:SalesRegion
          }
        }
      }
      layout row {
        tile company {
          value: "ID: " + ToText(SFDCAccounts:id)
        }
      }
      layout row {
        tile company {
          value: "Earliest Renewal Date: " + Left(ToText(SFDCAccounts:AccountRenewalDate), 10)
        }
      }
      layout row {
        tile company {
          value: "Renewals: " + SFDCAccounts:Agreement_Last_Dates
        }
      }
      // layout row {
      //   tile company {
      //     value: "On-Premise Renewal: " + ToText(CalendarDate(SFDCAccounts:AccountRenewalDateOnPremise))
      //   }
      //}
    }
  }
  widget summary {

    infobox {
      label: "Overall Risk Summary"
      info: "The top level summary widget provides a quick view of the current performance within the dimensions used to identify level of risk for the selected account. The Risk calculation is a weighted index that examines the customer's feelings (as measured by our Empower program), behavior (measured through our financial and Salesforce data), and our alignment with their feelings (as measured by our VoCe program)."
    }

    size: large
    table: SFDCAccounts:

    tile risk {
      label: "Overall Risk"
      showThermometer: false
      value: SFDCAccounts:overallIndex
      textValue: SFDCAccounts:overallHealthRiskCategory
      min: 0
      max: 10
      target: @targets.indexScore
      //renewal: SFDCAccounts:AccountRenewalDate
      revenue: SFDCAccounts:ltrL12MRev
      revenueLabel: "Last 12 mnths Rev"

    }
    tile metric {
      label: "Client Behaviour"
      value: SFDCAccounts:clientBehaviourIndex
      target: @targets.indexScore
    }
    tile metric {
      label: "Client Feeling"
      value: SFDCAccounts:clientFeelingIndex
      target: @targets.indexScore
    }

    tile metric {
      label: "Team Feeling"
      value: SFDCAccounts:teamFeelingIndex
      target: @targets.indexScore
    }
    tile casesStatus {
      open: count(cases:CaseId)
      overdue: count(cases:overdue, cases:overdue = "Yes")
    }
    tile casesStatus {
      label: "Open Support tickets"
      open: sum(TicketSummary:count, TicketSummary:StatusId = 1)
      overdue: sum(TicketSummary:count, TicketSummary:StatusId = 1)
      showOverdueText: false

    }
  }

  widget contactList {
    label: "Account Contacts: Latest Response"
    infobox {
      label: "Account Contacts: Latest Response"
      info: "The Contacts widget provides a list of all contacts currently associated with this account within Salesforce."
    }

    view metric #npsgroup {
      backgroundColorFormatter: backgroundColorFormatterNPSgroup
      valueColorFormatter: valueColorFormatterNPSgroup
    }

    table: contacts:
    sortColumn: lastResponse
    sortOrder: descending
    size: large
    navigateTo: "Contact Overview"

    column value #name {
      label: "Name"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }
    // column value #country {
    //   label: "Country"
    //   value: contacts:MailingCountry
    // }
    column date #lastResponse {
      label: "Last Feedback Date"
      value: last(relationship:interview_start, relationship:interview_start, _IsNull(relationship:Q1) = false)
      align: center
    }
    column metric #nps {
      label: "NPS Group"
      value: IIF(last(score(relationship:Q1), relationship:interview_start, _IsNull(relationship:Q1) = false) >= 0, last(score(relationship:Q1), relationship:interview_start, _IsNull(relationship:Q1) = false), -1)
      align: center
      view: npsgroup
      target: 9
      format: NPSgroupsContacts
    }
    column date #lastInvited {
      label: "Last Invite Date"
      value: last(respondent:smtpStatusDate, respondent:smtpStatusDate)
      align: center
    }
    column value #comments {
      label: "Recent Comment"
      value: last(relationship:Q2, relationship:interview_start, _IsNull(relationship:Q1) = false)
    }

    column value #noCases {
      label: "Total Cases"
      value: count(cases:CaseId)
      align: center
    }

    column value #overdueCases {
      label: "Overdue Cases"
      value: count(cases:CaseId, cases:overdue = "Yes")
      align: center
    }

  }

  widget dataGridBeta #clientBehaviourSummary2 {
    label: "Client Behaviour (Last 12 months)"
    size: large

    // suppressRule {
    //   criteria: COUNT(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRel) = 0
    //   label: "No responses to the relationship survey in the last 12 months"
    // }

    infobox {
      label: "Client Behaviour"
      info: "The Client Behaviour widget provides a view of all of the operational level data used to determine the overall Client Behavior score.

**Client Behavior**

- Spend Trend = Change in revenue in last 12 months
- Product Usage = RVA's used compared to those sold
- Response Rate = For Relationship survey only,
- Marketing Engagement = Index based on data available in SFDC
    - **Usage does not include usage of RVAs for Active Dashboards**"
    }

    view comparativeStatistic #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
    }

    view comparativeStatistic #adoptionlevelbehaviour {
      backgroundColorFormatter: adoptionTextBgColorFormatter
      valueColorFormatter: adoptionTextColorFormatter
    }

    view comparativeStatistic #index {
      backgroundColorFormatter: backgroundColorFormatterIndex
      valueColorFormatter: valueColorFormatterIndex
    }

    row {
      //label: "Client Feeling"

    }
    column {
      label: "Client Behav."
      cell {
        value: iif(SFDCAccounts:clientBehaviourIndex >= 0, SFDCAccounts:clientBehaviourIndex, -1)
        target: 8
        view: index
      }
    }
    column {
      label: "User Adopt."
      cell {
        value: IIF(@index.UserAdoption >= 0, @index.UserAdoption, -1)
        format: usertrend
        view: adoptionlevelbehaviour
        target: 10
      }
    }
    column {
      label: "RVA used / purch."
      cell {
        value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)"))
      }
    }
    column {
      label: "Mrkt Eng."
      cell {
        value: @index.LeadScore
        format: LeadScore
        view: adoptionlevelbehaviour
        target: 10
      }

    }
    column {
      label: "# Mrkt Contacts"
      cell {
        value: count(SFDCMarketLeads:Id)
        format: nodecimal
        align: center
      }
    }
    column {
      label: "Response Rate"
      cell {
        value: SFDCAccounts:responseRateL12M
        format: percentage
        align: center
      }
    }
    column {
      label: "Spend Trend"
      cell {
        value: @index.SpendTrend
        format: spendtrend
        view: adoptionlevelbehaviour
        target: 10
      }
    }
    column {
      label: "Rev. Diff (%)"
      cell {
        value: SFDCAccounts:revDiff
        //format: percentageonedecimal
        align: right
      }
    }

    column {
      label: "Last 12Mth Rev."
      cell {
        value: SFDCAccounts:ltrL12MRev
        format: UScurrency
        align: right
      }
    }
    column {
      label: "Prev 12Mth Rev."
      cell {
        value: SFDCAccounts:ltrP12MRev
        format: UScurrency
        align: right
      }
    }
    column {
      label: "Future - Best Case / Closed / Commit / Pipeline"
      cell {
        value: SFDCAccounts:FutureBCCCP
        format: UScurrency
        align: right
      }
    }

  }

  widget dataGridBeta #clientFeelingSummary2 {
    label: "Client feeling (Last 12 months average)"
    size: medium

    // suppressRule {
    //   criteria: COUNT(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRel) = 0
    //   label: "No responses to the relationship survey in the last 12 months"
    // }

    infobox {
      label: "Client Feeling"
      info: "The Client Feeling widget provides a consolidated view of the survey questions/responses from the Client Relationship and Implementation surveys that are currently being used to determine the Client Feeling score.

**Currently measured by Relationship Survey only**
- NPS (5%)
- Fulfils my Needs (40%)
- Delivers value to my organisation (15%)
- Satisfaction with the team (10%)
- Satisfaction with the technology (30%)
 *We will incorporate Implementation, Support & Training surveys into this metric*"
    }

    view comparativeStatistic #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
    }

    view comparativeStatistic #index {
      backgroundColorFormatter: backgroundColorFormatterIndex
      valueColorFormatter: valueColorFormatterIndex
      fontsize: large
    }

    row {
      //label: "Client Feeling"
    }

    column {
      label: "Client Feeling"
      cell {
        value: iif(SFDCAccounts:clientFeelingIndex >= 0, SFDCAccounts:clientFeelingIndex, -1)
        target: 8
        view: index
      }
    }
    column {
      label: "# Responses"
      cell {
        value: COUNT(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.L12MonthRel)
        format: integerDefaultFormatter
      }
    }
    column {
      label: "Likelihood to recommend"
      cell {
        value: iif(SFDCAccounts:NPSavg >= 0, SFDCAccounts:NPSavg, -1)
        target: 9
        view: metric
      }

    }
    column {
      label: "Support Business Needs"
      cell {
        value: iif(SFDCAccounts:NEEDSavg >= 0, SFDCAccounts:NEEDSavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Added Value"
      cell {
        value: iif(SFDCAccounts:VALUEavg >= 0, SFDCAccounts:VALUEavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Relationship Satisfaction"
      cell {
        value: iif(SFDCAccounts:RELavg >= 0, SFDCAccounts:RELavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Technology Satisfaction"
      cell {
        value: iif(SFDCAccounts:TECHavg >= 0, SFDCAccounts:TECHavg, -1)
        target: 9
        view: metric
      }
    }
  }

  widget dataGridBeta #teamFeelingSummary2 {

    // suppressRule {
    //   criteria: count(teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC) = 0
    //   label: "No responses to the team check survey in the last 12 months"
    // }

    infobox {
      label: "Team Feeling"
      info: "The Team Feeling widget provides a consolidated view of the survey questions/responses from the latest internal Health Check (and Implementation surveys - TBC) used to determine the Team Feeling score.

**Team Feeling**

*Currently measured by Account Manager perception of *

- NPS (5%)
- Liklihood to renew (40%)
- Recognise benefits across the organisation (15%)
- Confirmit support experience (40%)"
    }

    label: "Team feeling (Latest response in last 12 months)"
    size: medium

    view comparativeStatistic #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small

    }
    view comparativeStatistic #index {
      backgroundColorFormatter: backgroundColorFormatterIndex
      valueColorFormatter: valueColorFormatterIndex
    }
    row {
      //label: "Client Feeling"

    }
    column {
      label: "Team Feeling"
      cell {
        value: iif(SFDCAccounts:teamFeelingIndex >= 0, SFDCAccounts:teamFeelingIndex, -1)
        target: 8
        view: index
      }
    }
    column {
      label: "Latest Response Received (L12 Months)"
      cell {
        value: last(teamcheck:interview_start, teamcheck:interview_start, _IsNull(teamcheck:Q1) = false AND @daterange.L12MonthTC)
        format: dateDefaultFormatter

      }
    }
    column {
      label: "Likelihood to recommend"
      cell {
        value: iif(SFDCAccounts:tNPSavg >= 0, SFDCAccounts:tNPSavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Likelihood To Renew"
      cell {
        value: iif(SFDCAccounts:RENEWavg >= 0, SFDCAccounts:RENEWavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Recognises benefits"
      cell {
        value: iif(SFDCAccounts:BENavg >= 0, SFDCAccounts:BENavg, -1)
        target: 9
        view: metric
      }
    }
    column {
      label: "Confirmit support experience"
      cell {
        value: iif(SFDCAccounts:EXPavg >= 0, SFDCAccounts:EXPavg, -1)
        target: 9
        view: metric
      }
    }

  }


  widget contactList {

    infobox {
      label: "Team Checks"
      info: "TBC."
    }

    label: "Team Check: History"

    table: teamcheck:
    sortColumn: lastResponse
    sortOrder: descending
    size: large

    navigateTo: TeamCheckResponse


    view metric #metric {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
    }

    view metric #npsgroup {
      backgroundColorFormatter: backgroundColorFormatterNPSgroup
      valueColorFormatter: valueColorFormatterNPSgroup
    }

    column value #name {
      label: "Name"
      value: teamcheck:AccountOwner
    }

    column date #lastInvited {
      label: "Invite Date"
      value: teamcheck:FirstMailedDate
      align: center
    }

    column date #lastResponse {
      label: "Feedback Date"
      value: teamcheck:interview_start
      align: center
    }
    column metric #nps {
      label: "NPS Group"
      value: score(teamcheck:Q1)
      view: npsgroup
      target: 9
      align: center
      format: NPSgroupsContacts
    }

    column metric #ltr {
      label: "Recommend"
      value: score(teamcheck:Q1)
      align: center
      target: 9
      view: metric
    }

    column metric #renew {
      label: "Renew"
      value: score(teamcheck:Q2)
      align: center
      target: 9
      view: metric
    }

    column metric #recognise {
      label: "Benefits"
      value: score(teamcheck:Q8)
      align: center
      target: 9
      view: metric
    }

    column metric #supportexerience {
      label: "Support"
      value: score(teamcheck:Q9)
      align: center
      target: 9
      view: metric
    }
  }

  widget dataGridBeta #Opportunities1 {
    label: "Last 24 Months Rolling & Future Opportunities"
    size: large

    filter expression {
      value: (Between(SFDCClosedOpportunities:CloseDate, AddYear(GetDate(), -2), GetDate()) AND SFDCClosedOpportunities:IsClosed = "true") OR SFDCClosedOpportunities:CloseDate > GetDate()
    }

    row cut {
      value: SFDCClosedOpportunities:Name + " (" + SFDCClosedOpportunities:Id + ")"
      total: none

    }

    column {
      label: "Opportunity Closed Date"

      cell {

        value: Max(SFDCClosedOpportunities:CloseDate)
        format: dateDefaultFormatter
      }
    }
    column {
      label: "Opportunity Status"

      cell {
        value: Max(SFDCClosedOpportunities:ForecastCategoryName)
      }
    }
    column {
      label: "Opportunity Amount ($)"
      cell {
        value: Sum(SFDCClosedOpportunities:Amount_USD)
        format: UScurrency
      }
    }
  }

  widget chart #eJournalTicketCategories2 {
    label: "Support Tickets by Category (last 12 months)"
    size: large
    legend: topCenter
    layout: vertical
    scroll: auto
    chart bar {
      mode: stacked
      dataLabel: valueThenPercent
    }
    series {
      value: sum(TicketSummary:count)
      breakdownBy cut {
        value: IIF(TicketSummary:StatusId = 2, "Closed Tickets", "Open Tickets")
      }
    }
    category cut #categoryName {
      value: TicketCategories:fullname
      label: "Ticket Categories"
    }
    axis category {
      //orientation: 90
    }

    margin {
      left: 200
    }
    axis primary {
    //  axisLine: false

    }
  }
  widget markdown {
    label: " "
    markdown: "- Please note that the initial mapping of SFDC Acounts to Horizons accounts were done manually so there may be a small % of accounts that are unmapped or mapped incorrectly.
    - Only On-Demand usage data is currently included.
    - Additionally the usage data e.g. number RVAs used vs purchased, is not complete because usage data is not available for all products in Horizons, only Reportal and Dashboard / Instant Analytics is covered in the results."

    size: large
  }

  widget contactSurveyResponse {
    label: "Horizons Information"
    size: large
    table: SFDCAccounts:

//     summary {
//       rows: 5

//       tile list #list1 {
//         item value {
//           value: SFDCAccounts:Id
//           label: "Account ID"
//         }
//         item value {
//           value: SFDCAccounts:AccountOwnerName
//           label: "Account Owner"
//         }
//         item date {
//           label: "Account Renewal Date"
//           value: SFDCAccounts:AccountRenewalDate
//           format: dateDefaultFormatter
//         }
//       }
//       tile list #list2 {
//         item value {
//           value: SFDCAccounts:SalesRegion
//           label: "Region"
//         }
//         item value {
//           value: SFDCAccounts:ltrL12MRev
//           format: UScurrency
//           label: "Revenue Last 12 Months"
//         }
//         item value {
//           value: SFDCAccounts:ltrP12MRev
//           format: UScurrency
//           label: "Revenue Previous 12 Months"
//         }
//       }
//     }
//  // end of summary

    tab {
      label: "SITES SUMMARY"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Sites"
          value: ToText("EURO:" + IIF(count(usageAccounts:Id, usageAccounts:site = "euro") > 0, "YES", "No") + " / US:" + IIF(count(usageAccounts:Id, usageAccounts:site = "us") > 0, "YES", "No") + " / AUS:" + IIF(count(usageAccounts:Id, usageAccounts:site = "aus") > 0, "YES", "No") + " /CA:" + IIF(count(usageAccounts:Id, usageAccounts:site = "ca") > 0, "YES", "No") + " / HK:" + IIF(count(usageAccounts:Id, usageAccounts:site = "hk") > 0, "YES", "No"))
        }
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id)
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize)
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize)
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData)
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData)
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData)
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate())
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate())
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52) > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51) > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56) > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3) > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55) > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20) > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37) > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49) > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63) > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34) > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61) > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57) > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39) > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44) > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25) > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62) > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54) > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28) > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53) > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21) > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7) > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29) > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64) > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8) > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27) > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33) > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16) > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40) > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48) > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24) > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2) > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46) > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60) > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59) > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58) > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45) > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50) > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22) > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22) > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives") > 0, "YES", "No")
        }

      }

    }

    tab {
      label: "EUROPE"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "euro")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "euro")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "euro")
          format: nodecimal
        }

        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "euro")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "euro")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "euro")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "euro"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "euro")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "euro")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "euro") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "USA"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "us")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "us")
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "us")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "us")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "us")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "us"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "us")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "us")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "us") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "us") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "AUSTRALIA"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "aus")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "aus")
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "aus")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "aus")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "aus")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "aus"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "aus")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "aus")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "aus") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "CANADA"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "ca")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "ca")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "ca")
          format: nodecimal
        }

        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "ca")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "ca")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "ca")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "ca")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "ca") > 0, "YES", "No")
        }
      }
    }

    tab {
      label: "HONG KONG"
      tile list {
        label: "Licenses & Storage"
        item comment {
          label: "# Horizons Companies"
          value: count(usageAccounts:Id, usageAccounts:site = "hk")
        }
        item comment {
          label: "File Libary Used Size"
          value: sum(usageAccountStatistics:FileLibraryUsedSize, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "File Libary Limit"
          value: sum(usageAccountStatistics:FileLibraryLimitSize, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "Smart Hub Data"
          value: sum(usageAccountStatistics:SmartHubData, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "Survey Data"
          value: sum(usageAccountStatistics:SurveyData, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "Multimedia Data"
          value: sum(usageAccountStatistics:MultimediaData, usageAccounts:site = "hk")
          format: nodecimal
        }
        item comment {
          label: "# Professional Users"
          value: count(usageProfessionalUsers:Id, usageProfessionalUsers:DateExpires > GetDate() AND usageAccounts:site = "hk")
        }
        item comment {
          label: "# Translator Users"
          value: count(usageTranslatorUsers:Id, usageTranslatorUsers:DateExpires > GetDate() AND usageAccounts:site = "hk")
        }
        item comment {
          label: "# RVA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "hk")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report View Access (RVA)" AND usageAccounts:site = "hk"))
        }
        item comment {
          label: "# RAA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "hk")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Analyst Access (RAA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# RDA used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "hk")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Report Design Access (RDA)" AND usageAccounts:site = "ca"))
        }
        item comment {
          label: "# Dashboard/Instant Analytics licenses used vs purchased"
          value: ToText(sum(usageReportalLicenses:Users, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "ca")) + " / " + ToText(sum(usageReportalLicenses:Purchased, usageReportalLicenses:Type = "Dashboard/Instant Analytics" AND usageAccounts:site = "hk"))
        }
        item comment {
          label: "CATI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CATI Seats" AND usageAccounts:site = "hk")
        }
        item comment {
          label: "CAPI Seats"
          value: sum(usageLicenses:Users, usageLicenses:Type = "CAPI Seats" AND usageAccounts:site = "hk")
        }
      }
      tile list {
        label: "Enabled Features"
        item comment {
          label: "Actions"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 52 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Active Dashboards"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 51 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "AskMe Offline Survey Completion App"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 56 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Basic Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 3 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Business User Access to Hierarchy Management"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 55 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CAPI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 20 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CATI"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 37 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CATI Call Centers"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 49 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CATI IVR"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 63 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Concurrent Sampling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 34 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for MS Dynamics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 61 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connector for Salesforce"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 57 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Data Processing"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 39 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Database Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 44 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Dedicated IP"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 25 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Digital Feedback"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 62 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Discovery Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 54 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "DomainKeys"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 28 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Feature Toggling"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 53 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "File Library"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 21 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "FTP for file transfer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 7 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Kiosk"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 29 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Native Survey SDK"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 64 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "PGP Encryption"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 8 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Professional Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 27 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Questionnaire Reviewer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 33 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Random Data Generator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 16 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Sample Only"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 40 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Short Url"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 48 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Single Sign On"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 24 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Spell checker"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 2 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Standard Panel"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 46 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for B2B Account Health"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 60 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Deployment for Employee Pulse"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 59 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Studio Designer"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 58 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Survey Router"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 45 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Text Analytics"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 50 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Transaction Types"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Translator"
          value: IIF(count(usageActivatedModules:, usageActivatedModules:ModuleId = 22 AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
      }
      tile list {
        label: "Flex Extensions"
        item comment {
          label: "Android Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Android Surveys" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Confirmit Question Extensions"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Confirmit Question Extensions" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "CRM Connect for SalesForce"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "CRM Connect for SalesForce" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Email Frequency Filter"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Email Frequency Filter" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "E-mail Opt Out"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "E-mail Opt Out" OR usageFlexExtensions:Name = "Email Opt Out") AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "FRend"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "FRend" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Geolocation"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Geolocation" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "iPhone Surveys"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "iPhone Surveys" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Language Translator"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Language Translator" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Mobile Portal"
          value: IIF(count(usageFlexExtensions:, ((usageFlexExtensions:Name = "Mobile Portal Prototype" OR usageFlexExtensions:Name = "MobilePortal") OR usageFlexExtensions:Name = "MobilPortal") AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "SMS Surveys"
          value: IIF(count(usageFlexExtensions:, (usageFlexExtensions:Name = "SMS Surveys" OR usageFlexExtensions:Name = "SmsSurveys") AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Social Data Import"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Social Data Import" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "SurveyBuddy"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "SurveyBuddy" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Translation Review"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Translation Review" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "TRC Speeder"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TRC Speeder" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "TrueSample"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "TrueSample" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Ugam ENRAPTURE"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Ugam ENRAPTURE" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
        item comment {
          label: "Virtual Incentives"
          value: IIF(count(usageFlexExtensions:, usageFlexExtensions:Name = "Virtual Incentives" AND usageAccounts:site = "hk") > 0, "YES", "No")
        }
      }
    }

  }
}

page account #TeamCheckResponse {
  modal: true

  label: "Team Check Response"

  widget contactSurveyResponse {
    view title #defaultSurveyResponseTitle {
    }
    size: medium


    surveyResponseTitle {
      tile title #rt {
        value: SFDCAccounts:AccountOwnerName + " - Team Check Survey"
        surveyName: "Team Check Survey"
        view: defaultSurveyResponseTitle
      }
    }

    summary {
      rows: 4
      tile list #list1 {
        item value {
          value: teamcheck:status
          label: "Status"
        }
        item date {
          value: teamcheck:interview_start
          label: "Feedback Received"
          format: long
        }
      }
      tile list #list2 {
        item value {
          value: "Team Check Survey"
          label: "Source"
        }
        item value {
          value: teamcheck:responseid
          label: "Response ID"
        }
      }
    }
 // end of summary

    tab {
      label: "Responses"
      tile list {
        label: " "
        item comment {
          label: "Region"
          value: SFDCAccounts:SalesGroupRegion
        }
        item comment {
          label: "Team"
          value: SFDCAccounts:SalesRegion
        }
        item comment {
          label: "Company name"
          value: SFDCAccounts:Name
        }
        item comment {
          label: "Customer Type"
          value: SFDCAccounts:ClientType
        }
        item comment {
          label: "Industry"
          value: SFDCAccounts:Industry
        }
      }
      tile list {
        label: "Survey Responses"
        item bar {
          label: "Likelihood to Recommend"
          value: score(teamcheck:Q1)
        }
        item bar {
          label: "Likelihood to Renew"
          value: score(teamcheck:Q2)
        }
        item comment {
          label: "Why not renew?"
          value: teamcheck:Q3
        }
        item comment {
          label: "How to keep?"
          value: teamcheck:Q4
        }
        item bar {
          label: "Spend Potential"
          value: score(teamcheck:Q5)
        }
        item comment {
          label: "Increase Spend?"
          value: teamcheck:Q6
        }
        item comment {
          label: "Decrease Spend?"
          value: teamcheck:Q7
        }
        item bar {
          label: "Recognise Benefits"
          value: score(teamcheck:Q8)
        }
        item bar {
          label: "Support Experience"
          value: score(teamcheck:Q9)
        }
        item comment {
          label: "Support Experience comments"
          value: teamcheck:Q10
        }
        item bar {
          label: "Dependency on Services"
          value: score(teamcheck:Q11)
        }
        item bar {
          label: "Dependency on Support"
          value: score(teamcheck:Q12B)
        }
      }
    }
  }
}

page contact #ContactOverview {
  label: "Contact Overview"

  modal: true

  widget title {
    table: contacts:
    view icon #icon {
      size: "60"
      roundedCorner: true
    }

    layout column {
      tile value #logo {
        value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/magdalenas/defaultLogo.PNG"//"http://is1.mzstatic.com/image/thumb/Purple71/v4/89/51/f4/8951f4f1-fd6b-fa59-38b2-191140473b9a/source/175x175bb.jpg"
        view: icon
      }
    }
    layout column {
      layout row {
        tile value #firstName {
          value: contacts:FirstName
        }
        tile value #lastName {
          value: contacts:LastName
        }
        tile role {
          value: contacts:ContactRole
        }
      }
      layout row {
        tile company {
          value: SFDCAccounts:Name
          navigateTo: "Account Overview"
        }
      }
    }
  }

  widget summary {

    infobox {
      label: "Contact Summary"
      info: "The Contact Summary widget provides a window into some of the information captured for this contact within Salesforce, along with some key metrics associated with the overall risk calculation for the account (likelihood to renew, response rate). The email link is live, and allows you to email the contact directly from this screen."
    }

    size: large
    table: contacts:
    tile contactDetails #cc {
      title: contacts:Title
      role: contacts:ContactRole
      email: contacts:email
      phone: contacts:Phone
      industry: contacts:Industry
    }

    tile accountDetails #cc4 {
      accountOwner: SFDCAccounts:AccountOwnerName
      region: contacts:WorldRegion
      revenue: SFDCAccounts:ltrL12MRev
      renewalDate: SFDCAccounts:AccountRenewalDate

    }

    tile metric #a {
      label: "LTR"
      value: round(average(score(relationship:Q1)), 1)
      target: 9
    }

    tile responseRate {
      label: "Response Status"
      invites: COUNT(respondent:respid, @filter.isSent)
      responses: COUNT(relationship:responseId, @filter.isPartial OR @filter.isResponded)
    }

    tile casesStatus {
      label: Cases
      open: count(cases:CaseId)
      overdue: 0
    }
  }

  widget contactSurveys {

    infobox {
      label: "Feedback History"
      info: "The Feedback History widget lists all feedback responses captured for this contact from {what time frame?}. This is valuable in understanding how/if a specific contact's perception has shifted over time. The blue "
      Resend #linkprovidestheAccountManagerwiththeabilitytoresendasurveyiftheoriginalsurveywasntreceivedbythecustomerorifanadditionalreminderisrequired
    }

    label: "Feedback History"
    table: respondent:
    sortColumn: surveyDate
    sortOrder: descending
    size: medium
    navigateTo: "Response"

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    // column value #respondent {
    //   label: "Respid"
    //   value: respondent:respid
    // }
    // column value #lastRespidContact {
    //   label: "Last Resp ID Contact"
    //   value: contacts:LastRespondentId
    // }
    column date #inviteDate {
      label: "Request Date"
      value: respondent:FirstEmailedDate
      format: dateDefaultFormatter
    }
    column date #surveyDate {
      label: "Response Date"
      value: relationship:interview_start
      format: dateDefaultFormatter
    }

    column value #survey {
      label: "Survey"
      value: "Relationship"
    }
    column value #status {
      label: "Status"
      value: respondent:responseStatus
    }

    column link #Resend {
      label: "Resend invite"
      value: IIF(relationship:status = "incomplete" OR _IsNull(relationship:status), IIF(respondent:respid = Last(respondent:respid, respondent:respid) AND @daterange.L3MonthRelResp, "Resend", ""), "")
      link surveyBlock #myLink {
        survey: p1850259384
        blockId: "Resend Invite"
        respid: respondent:respid
      }
    }

    column metric #ltr {
      label: "LTR"
      value: score(relationship:Q1)
      view: metrics
      target: 9
      align: center
    }

    column value #comments {
      label: "Comments"
      value: relationship:Q2
    }

  }

  widget accountCases {

    infobox {
      label: "Case History"
      info: "The Case History widget provides a list of all cases opened as a result of direct feedback from this contact from {what time frame?}"
    }

    label: "Case History"
    table: cases:
    size: medium
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #dateCreated {
      label: "Created"
      value: cases:DateCreated
      format: long
      align: center
    }
    column value #dateDue {
      label: "Due"
      value: cases:DateDue
      format: long
      align: center
    }

    column value #caseStatus {
      label: "Status"
      value: cases:lk_1545
    }
    column value #issuetype {
      label: "Issues Identified"
      value: cases:lk_1547
    }
    column value #link {
      label: "Action"
      value: cases:CaseLink
      view: link1
    }
  }

}

page #CustomerAlerts {
  label: "Customer Alerts"

  modal: true

  filter expression {
    value: @daterange.currentPeriodCases
    filtertype: "preAggregate"
  }

  widget barChart {


    infobox {
      label: "Issues Triggering Customer Alerts"
      info: "The Issues Triggering Customer Alerts widget highlights the status of all negative alerts stemming from the Relationship Survey and the Implementation survey from the last 12 months."
    }
    table: cases:
    label: "Issues Triggering Customer Alerts"
    size: large
    value: count(cases:caseId)
    //palette: "#0F5E7D","#FFBB5C","#CF2740","#ED4F34","#CCCCCC","#333333","#F58533"
    navigateTo: "Cases"
    category cut {
      value: cases:lk_1547
      removeEmpty: true
    }
    series cut {
      value: cases:lk_1545
    }
  }

  widget accountCases {

    infobox {
      label: "Cases"
      info: "The Cases widget provides a list of all cases from the Relationship survey and the Implementation survey, along with current status. Click on the blue ''View case' link to view the fully recorded details regarding that particular case."
    }

    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #accountName {
      label: "Account"
      value: SFDCAccounts:Name
    }

    column value #Contact {
      label: "Contact"
      value: contacts:FirstName + " " + contacts:LastName
    }

    column value #dateCreated {
      label: "Created"
      value: cases:DateCreated
      format: long
      align: center
    }
    column value #dateDue {
      label: "Due"
      value: cases:DateDue
      format: long
      align: center
    }
    column value #workflow {
      label: "Workflow"
      value: cases:Workflow
    }
    column value #caseStatus {
      label: "Status"
      value: cases:lk_1545
    }
    column value #issuetype {
      label: "Issues Identified"
      value: cases:lk_1547
    }
    column value #link {
      label: "Action"
      value: cases:CaseLink
      view: link1
    }
  }

}


page #Cases {
  label: "Cases"


  filter expression {
    value: @daterange.currentPeriodCases
    filtertype: "preAggregate"
  }

  modal: true

  widget accountCases {
    infobox {
      label: "Cases"
      info: "NA"
    }

    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #accountName {
      label: "Account"
      value: SFDCAccounts:Name
    }

    column value #Contact {
      label: "Contact"
      value: contacts:FirstName + " " + contacts:LastName
    }

    column value #dateCreated {
      label: "Created"
      value: cases:DateCreated
      format: long
      align: center
    }
    column value #dateDue {
      label: "Due"
      value: cases:DateDue
      format: long
      align: center
    }
    column value #workflow {
      label: "Workflow"
      value: cases:Workflow
    }
    column value #caseStatus {
      label: "Status"
      value: cases:lk_1545
    }
    column value #issuetype {
      label: "Issues Identified"
      value: cases:lk_1547
    }
    column value #link {
      label: "Action"
      value: cases:CaseLink
      view: link1
    }
  }

}

page #ResponseManagement {
  label: "Response Management"


  widget accountList {

    infobox {
      label: "Account Response Status"
      info: "The Account Response Status widget provides a list of accounts for whom surveys have been sent, with low response rate (less than 25% in the last 12 months). The lack of response/engagement could be an indicator of risk. Account Managers should pay close attention to any customers who are not providing at least one response to the Empower relationship survey during the year."
    }

    label: "Account Response Status"
    size: large
    table: SFDCAccounts:
    sortColumn: account
    sortOrder: ascending
    navigateTo: "Non Responders"

    take: 100
    paginationType: paging
    rowsPerPage: 100,150,200,250
    headerNumberOfLines: 4

    column value #account {
      label: "Account"
      value: SFDCAccounts:Name
      enableColumnFilter: true
    }
    column value #active {
      label: "Is Active"
      value: IIF(SFDCAccounts:ActiveClient = "True", "Yes", "No")
    }
    column value #accountrenewaldate {
      label: "Renewal Date"
      value: SFDCAccounts:AccountRenewalDate
      format: dateDefaultFormatter
    }
    column value #responseRateL12M {
      label: "Response Rate L12 months"
      value: SFDCAccounts:responseRateL12M
      format: percentage
    }
    column value #LastInvite {
      label: "Last Invite Sent"
      value: max(respondent:smtpStatusDate, @filter.isSent)
      format: dateDefaultFormatter
      align: center
    }
    column value #LastResponse {
      label: "Last Response"
      value: max(relationship:interview_start, @filter.isSent)
      format: dateDefaultFormatter
      align: center
    }
    column value #LastTeamCheck {
      label: "Last Team Check"
      value: max(teamcheck:interview_start, _IsNull(teamcheck:Q1) = false)
      format: dateDefaultFormatter
      align: center
    }
    column value #invites {
      label: "Total Invites"
      value: COUNT(respondent:respid, @filter.isSent)

    }
    column value #responses {
      label: "Total Responses"
      value: COUNT(relationship:responseId, @filter.isPartial OR @filter.isResponded)
    }
  }
}


page #AccountAlerts {

  filter expression {
    value: @daterange.currentPeriodCases
    filtertype: "preAggregate"
  }
  label: "Customer Alerts"
  widget barChart {


    infobox {
      label: "Issues Triggering Customer Alerts"
      info: "The Issues Triggering Customer Alerts widget highlights the status of all negative alerts stemming from the Relationship Survey and the Implementation survey from the last 12 months."
    }
    table: cases:
    label: "Issues Triggering Customer Alerts"
    size: large
    value: count(cases:caseId)
    palette: "#0F5E7D","#FFBB5C","#CF2740","#ED4F34","#CCCCCC","#333333","#F58533"
    navigateTo: "Cases"
    category cut {
      value: cases:lk_1547
      removeEmpty: true
    }
    series cut {
      value: cases:lk_1545
    }
  }

  widget accountCases {

    infobox {
      label: "Cases"
      info: "The Cases widget provides a list of all cases from the Relationship survey and the Implementation survey, along with current status. Click on the blue ''View case' link to view the fully recorded details regarding that particular case."
    }

    label: "Cases"
    table: cases:
    size: large
    sortColumn: dateCreated
    sortOrder: descending

    view link #link1 {
      label: "View case"
    }

    column value #accountName {
      label: "Account"
      value: SFDCAccounts:Name
    }

    column value #Contact {
      label: "Contact"
      value: contacts:FirstName + " " + contacts:LastName
    }

    column value #dateCreated {
      label: "Created"
      value: cases:DateCreated
      format: long
      align: center
    }
    column value #dateDue {
      label: "Due"
      value: cases:DateDue
      format: long
      align: center
    }
    column value #workflow {
      label: "Workflow"
      value: cases:Workflow
    }
    column value #caseStatus {
      label: "Status"
      value: cases:lk_1545
    }
    column value #issuetype {
      label: "Issues Identified"
      value: cases:lk_1547
    }
    column value #link {
      label: "Action"
      value: cases:CaseLink
      view: link1
    }
  }

}

page #NonResponders {
  label: "Non Responders"

  modal: true


  widget contactSurveys {

    infobox {
      label: "Accounts: Invite History"
      info: "NA"
    }


    label: "Accounts: Invite History"
    table: respondent:
    navigateTo: "Response"
    sortColumn: inviteDate
    sortOrder: descending
    size: large

    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
      //roundCorners:true
    }
    column value #name {
      label: "Contact"
      value: contacts:FirstName + " " + contacts:LastName
    }
    column value #account {
      label: "Account"
      value: SFDCAccounts:Name
    }
    column value #role {
      label: "Role"
      value: contacts:ContactRole
    }
    column date #inviteDate {
      label: "Invite Date"
      value: respondent:smtpstatusDate
      format: dateDefaultFormatter
    }
    column value #status {
      label: "Response Status"
      value: relationship:status
    }
    column link #Resend {
      label: "Resend invite"
      value: IIF(relationship:status = "incomplete" OR _IsNull(relationship:status), IIF(respondent:respid = Last(respondent:respid, respondent:respid) AND @daterange.L3MonthRelResp, "Resend", ""), "")
      link surveyBlock #myLink {
        survey: p1850259384
        blockId: "Resend Invite"
        respid: respondent:respid
      }
    }
    column date #surveyDate {
      label: "Response Date"
      value: relationship:interview_start
      format: dateDefaultFormatter
    }
  }
}

page #BusinessOverview {

  label: "Business Health"

  widget markdown {
    size: large
    markdown: "Results for Net Sales Performance and Renewal Rate only includes financial data up to Q3 2019.
- Net Sales Performance and Renewal Rate results are always based on in the last 12 months rolling from the 1st of the current month.

**Note:**
*Any filtering applied via the Filter toolbar is not applied to these widgets.*"
  }


  widget kpi {

    infobox {
      label: "Net Sales Performance (Q3 '19)"
      info: "The Net Sales Performance widget is a quick view of current performance against our net sales metric target for last completed financial quarter. The black line within the arc represents the target. If the color is green the metric is at or above the acceptable range of the target score. If the color is yellow, the metric is within an x% margin lower than target. If the target is red, the current metric is outside of an acceptable range below the target and requires attention."
    }

    filter expression {
      value: InQuarter(finance:Month, -2, -2)
    }

    label: "Net Sales Performance (Q3 '19)"
    size: small
    tile kpi {
      label: "Quota Achievement"
      value: @calculate.salesperformance
      target: 100
      min: 0
      max: 100
      format: percentage
      targetFormat: percentage
      gaugeColorFormat: NetSalesGauge
      tile value {
        label: "New Clients"
        value: finance:Noofnewclients
    //format: nodecimal
      }
    }
  }


  widget chart {

    infobox {
      label: "Net Sales Performance vs Renewal Rate last 5 quarters"
      info: "The Net Sales Performance widget represents quarterly net sales figures as a percentage of expected quota for the last 5 quarters."
    }

    // filter expression {
    //   value: @daterange.currentPeriodFin
    // }

    label: "Net Sales Performance vs Renewal Rate last 5 quarters"
    palette: "#2B3E50","#DF691A","#54bc23"

    size: medium
    legend: bottomCenter
    gridLines: none

    chart line {
      //lineType: basis
      dotSize: 5
    }
    removeEmptyCategories: true

    series #ss1 {
      value: @calculate.salesperformance
      format: percentage
      label: "Net Sales Performance"
    }
    series #ss2 {
      value: Sum(finance:RevenueRenewalRate) * 100
      format: percentage
      label: "Renewal Rate"
    }


    series #ss3 {
      value: 100
      format: valueDefaultFormatter
      label: "target"
      chart line {
        lineType: linear
        dotSize: 0
      }
    }

    category date {
      value: finance:month
      breakdownBy: calendarQuarter
      label: "Date"
      start: "-6 quarters" // THIS MEEDS TO BE DYNAMIC
      end: "0 days"
      format: quarterlabel
    }

  }


  widget kpi {

    infobox {
      label: "Renewal Rate"
      info: "The Renewal Rate widget is a quick view of the current response rate for the Empower relationship survey for last completed financial quarter. The black line within the arc represents the target. If the color is green the metric is at or above the acceptable range of the target score. If the color is amber, the metric is within an x% margin lower than target. If the target is red, the current metric is outside of an acceptable range below the target and requires attention."
    }

    filter expression {
      value: InQuarter(finance:Month, -2, -2)
    }
    label: "Renewal Rate (Q3 '19)"
    size: small
    tile kpi {
      label: "Renewal Achievement"
      value: finance:RevenueRenewalRate * 100
      target: finance:RevenueRenewalRateTarget * 100
      min: 0
      max: 100
      format: percentage
      targetFormat: percentage
      gaugeColorFormat: RenewalRateGauge

    }
  }

  widget markdown {
    size: large
    markdown: "Results for the NPS Performance Trend is only available as a global total.
    **Note:** Any filtering applied via the Filter toolbar is not applied to these widgets.*"
  }

  widget kpi {
    infobox {
      label: "Client NPS"
      info: "The Client NPS widget is a quick view of the current NPS scores coming through the Empower relationship survey for {what time frame?}. The black line within the arc represents the target. If the color is green the metric is at or above the acceptable range of the target score. If the color is yellow, the metric is within an x% margin lower than target. If the target is red, the current metric is outside of an acceptable range below the target and requires attention."
    }
    suppressRule {
      criteria: count(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.currentPeriodRel) = 0
      label: "No responses found"
    }

    label: "Client NPS"
    size: small
    tile kpi {
      label: "NPS"
      value: NPS(relationship:Q1, @daterange.currentPeriodRel) * 100
      format: onedecimal
      min: -100
      max: 100
      target: 20
      targetFormat: onedecimal
      gaugeColorFormat: npsGauge
      showRange: true
      tile value {
        label: "Responses"
        value: count(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.currentPeriodRel)
      }
      tile value {
        label: "Yearly change"
        value: NPS(relationship:Q1, @daterange.L12MonthRel) * 100 - NPS(relationship:Q1, @daterange.P12MonthRel) * 100
        format: onedecimal

      }
      tile value {
        label: ""
        value: IIF(NPS(relationship:Q1, @daterange.L12MonthRel) * 100 > NPS(relationship:Q1, @daterange.P12MonthRel) * 100, "UP", "DOWN")

      }

    }
  }

  widget chart {
    infobox {
      label: "NPS Performance"
      info: "The NPS Performance widget provides a month by month comparison of NPS scores between the external customer relationship survey and the internal health check survey over the past 12 months. Actual scores for each month can be seen by hovering over the data points on the chart."
    }

    // filter expression {
    //   value: @daterange.currentPeriodTRCom
    // }
    //animation: true
    label: "NPS Performance"
    palette: "#2B3E50","#DF691A","#54bc23"
    size: medium
    legend: bottomCenter
    gridLines: none
    removeEmptyCategories: true

    chart line {
      //lineType: basis
      dotSize: 5
    }

    series #ss1 {
      value: NPS(clientandteam:Q1, clientandteam:combined_sourceid = "p1850259384") * 100
      format: onedecimal
      label: "Client NPS"
    }
    series #ss2 {
      value: NPS(clientandteam:Q1, clientandteam:combined_sourceid = "p1860215844") * 100
      format: onedecimal
      label: "Internal Team NPS"
    }
    series #ss3 {
      value: 20
      format: valueDefaultFormatter
      label: "target"
      chart line {
        lineType: linear
        dotSize: 0
      }
    }

    category overlappingDate {
      value: clientandteam:RelationshipSurveyDate
      breakdownBy: calendarMonth
      format: monthlabel
      start: "-12 months" // THIS MEEDS TO BE DYNAMIC
      end: "0 days"
      startShift: "-12 month"
      endShift: "0 month"

    }
  }


  widget kpi {

    infobox {
      label: "Internal Team NPS"
      info: "The Internal Team NPS widget is a quick view of the current NPS score as represented in Health Check surveys completed by the Account Managers for {what time frame?}. The black line within the arc represents the target. If the color is green the metric is at or above the acceptable range of the target score. If the color is yellow, the metric is within an x% margin lower than target. If the target is red, the current metric is outside of an acceptable range below the target and requires attention."
    }

    suppressRule {
      criteria: count(teamcheck:responseid, _IsNull(teamcheck:Q1) = false AND @daterange.currentPeriodTC) = 0
      label: "No responses found"
    }

    label: "Internal Team NPS"
    size: small
    tile kpi {
      label: "NPS"
      value: NPS(teamcheck:Q1, @daterange.currentPeriodTC) * 100
      format: onedecimal
      min: -100
      max: 100
      target: 20
      targetFormat: onedecimal
      showRange: true
      gaugeColorFormat: npsGauge
      tile value {
        label: "Responses"
        value: count(teamcheck:responseid, _IsNull(teamcheck:Q1) = false AND @daterange.currentPeriodTC)
      }
      tile value {
        label: "Yearly change"
        value: NPS(teamcheck:Q1, @daterange.L12MonthTC) * 100 - NPS(teamcheck:Q1, @daterange.P12MonthTC) * 100
        format: onedecimal
      }
      tile value {
        label: ""
        value: IIF(NPS(teamcheck:Q1, @daterange.L12MonthTC) * 100 > NPS(teamcheck:Q1, @daterange.P12MonthTC) * 100, "UP", "DOWN")
      }
    }
  }

  widget accountList {

    suppressRule {
      criteria: count(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.currentPeriodRel) + count(teamcheck:responseid, _IsNull(teamcheck:Q1) = false AND @daterange.currentPeriodTC) = 0
      label: "No responses found"
    }

    infobox {
      label: "How Are We Performing Across Regions"
      info: "The 'How Are We Performing Across Regions' widget represents current NPS scores {for what time period?} rolled up to the region level, with the ability to drill down through the regional account management hierarchy down to the account level."
    }

    label: "How Are We Performing Across Regions"
    table: hierarchy:
    hierarchy: hierarchy:21039

    size: large
   // sortColumn: hierarchy

    view metric #metriccell {
      backgroundColorFormatter: backgroundColorFormatterNPS
      valueColorFormatter: valueColorFormatterNPS
      //fontSize: large

    }

    column hierarchy {
      label: "Region"
      value: hierarchy:language_text
      removeEmpty: true
    }
    column metric {
      label: "Client NPS"
      value: NPS(relationship:Q1, @daterange.currentPeriodRel) * 100
      format: onedecimal
      target: @targets.NPS
      view: metriccell

    }
    column value {
      label: "# Responses"
      value: Count(relationship:Q1, @daterange.currentPeriodRel)
      format: onedecimal
    }
    column value {
      label: "Yearly change"
      value: NPS(relationship:Q1, @daterange.L12MonthRel) * 100 - NPS(relationship:Q1, @daterange.P12MonthRel) * 100
      format: onedecimal
    }

    column metric {
      label: "Internal Team NPS"
      value: NPS(teamcheck:Q1, @daterange.currentPeriodTC) * 100
      format: onedecimal
      target: @targets.tNPS
      view: metriccell
    }
    column value {
      label: "# Responses"
      value: Count(teamcheck:Q1, @daterange.currentPeriodTC)
      format: onedecimal
    }
    column value {
      label: "Yearly change"
      value: NPS(teamcheck:Q1, @daterange.L12MonthTC) * 100 - NPS(teamcheck:Q1, @daterange.P12MonthTC) * 100
      format: onedecimal
    }
  }

  widget markdown {
    size: large
    markdown: "Key metrics across the customer journey will be rolled into Empower in phases. Metrics listed below without data are scheduled for phases 2/3."
  }
  widget metricsBeta {

    infobox {
      label: "Research"
      info: "The Research widget highlights key metrics that inform on performance with our customers and prospects as they are researching and evaluating our offerings. *Does marketing have text describing their engagement score and the "
      Resend #linkprovidestheAccountManagerwiththeabilitytoresendasurveyiftheoriginalsurveywasntreceivedbythecustomerorifanadditionalreminderisrequired
    }

    view metricWithBar #metric {
      valueColorFormatter: acrossTheJourney
      showThermometer: false
    }

    view metricWithBar #metriccell {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      showThermometer: false
      fontSize: small
      roundCorners: false
    }

    label: "Research"
    size: small
    tile header {
      item title {
        value: "KPI"
        rowHeader: true
      }
      item title {
        value: "Average"
        rowHeader: true
      }
    }
    tile row {
      item value {
        value: "Marketing Engagement"
      }
      item metric {
        value: @index.LeadScore //average(LeadScore:mkto71_Lead_Score)
        view: metriccell
        target: 100
        format: LeadScore
      }
    }
    tile row {
      item value {
        value: "Confirmit.com Easy Score"
      }
      item metric {
        value: average(score(website:Q2.1))
        target: 8
        view: metriccell
      }
    }

    tile row {
      item value {
        value: "Funnel Progress"
      }
      item metric {
        value: ""
        view: metric
        target: 7
      }
    }
  }

  widget metricsBeta {

    infobox {
      label: "Decide"
      info: "The Decide widget highlights key metrics that inform on performance with our customers and prospects as they make their decision to proceed with, or decline to move forward with, our offerings. *Is there anything we can add regarding expected targets for SQL (and the other metrics)? Along with a short blurb about what is intended with this metric?  Metrics in green are in line with goals. Metrics in yellow are outside the range of being acceptable and should be monitored, but no action is required. Metrics in red are out of range of the expected goal and should be addressed."
    }

    view metricWithBar #metric {
      valueColorFormatter: acrossTheJourney
      showThermometer: false
    }

    view metricWithBar #metriccell {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      showThermometer: false
      fontSize: small
      roundCorners: false
    }

    label: "Decide"
    size: small
    tile header {
      item title {
        value: "KPI"
        rowHeader: true
      }
      item title {
        value: "Average"
        rowHeader: true
      }
    }
    tile row {
      item value {
        value: "Conversion Rate"
      }
      item metric {
        value: ""
        target: 100
        view: metric
      }
    }
    tile row {
      item value {
        value: "SQL Quota Achieved"
      }
      item metric {
        value: finance:SQLquotaachievement * 100
        view: metriccell
        target: 100
        format: percentage
      }
    }
    tile row {
      item value {
        value: "Revenue to Target"
      }
      item metric {
        value: ""
        view: metric
        target: 100
      }
    }
    tile row {
      item value {
        value: "Win/Loss Completion"
      }
      item metric {
        value: "" //average(score(relationship:Q9.1))
        view: metric
        target: 7
      }
    }
    tile row {
      item value {
        value: "New Accounts"
      }
      item metric {
        value: finance:Noofnewclients
        view: metriccell
        target: 7
      }
    }
  }

  widget metricsBeta {

    infobox {
      label: "Use"
      info: "The Use widget highlights key metrics that inform on performance with our customers and prospects as they are using our product and engaged with the teams that provide them with service. *How are we deriving user adoption? Is it based on usage somehow? The other 4 metrics are based on results from the implementation surveys provided to customers following an initial implementation or subsequent project. Metrics in green are in line with goals. Metrics in yellow are outside the range of being acceptable and should be monitored, but no action is required. Metrics in red are out of range of the expected goal and should be addressed."
    }

    view metricWithBar #metric {
      valueColorFormatter: acrossTheJourney
      showThermometer: false
    }
    view metricWithBar #metriccell {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      showThermometer: false
      fontSize: small
    }

    view metricWithBar #adoptionlevelbehaviour {
      backgroundColorFormatter: adoptionTextBgColorFormatter
      valueColorFormatter: adoptionTextColorFormatter
      showThermometer: false
    }

    label: "Use"
    size: small
    tile header {
      item title {
        value: "KPI"
        rowHeader: true
      }
      item title {
        value: "Average"
        rowHeader: true
      }
    }
    tile row {
      item value {
        value: "User Adoption"
      }
      item metric {
        value: IIF(average(@index.UserAdoption) >= 0, average(@index.UserAdoption), -1)
        format: usertrend
        view: adoptionlevelbehaviour
        target: 10
      }
    }

    // CANNOT DO THIS BECAUSE WE CANNOT ADD IMPLEMENTATION SOURCES.
    tile row {
      item value {
        value: "Implementation Met Needs"
      }
      item metric {
        value: ""// average(score(implementClient:C_Met_Needs.1))
        target: 8
        view: metriccell
      }
    }
    tile row {
      item value {
        value: "Relationship Satisfaction"
      }
      item metric {
        value: average(score(relationship:Q4), @daterange.currentPeriodRel)
        view: metriccell
        target: 8
      }
    }
    tile row {
      item value {
        value: "Technology Satisfaction"
      }
      item metric {
        value: average(score(relationship:Q7), @daterange.currentPeriodRel)
        view: metriccell
        target: 7
      }
    }
    tile row {
      item value {
        value: "Support Satisfaction"
      }
      item metric {
        value: ""
        view: metric
        target: 7
      }
    }
  }

  widget metricsBeta {

    infobox {
      label: "Renew"
      info: "The Renew widget highlights key metrics that inform on performance with our customers and prospects as they are considering whether or not to continue doing business with Confirmit. *Are renewal rate and growth rate YTD? Past 12 months? The likelihood to renew and supports needs metrics are derived from the current Empower relationship survey for {what time frame?}. Metrics in green are in line with goals. Metrics in yellow are outside the range of being acceptable and should be monitored, but no action is required. Metrics in red are out of range of the expected goal and should be addressed."
    }

   // viaStrategy: shortest

    table: SFDCAccounts:

    view metricWithBar #metric {
      valueColorFormatter: acrossTheJourney
      showThermometer: false
    }
    view metricWithBar #metriccell {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      showThermometer: false
      fontSize: small
    }
    label: "Renew"
    size: small
    tile header {
      item title {
        value: "KPI"
        rowHeader: true
      }
      item title {
        value: "Average"
        rowHeader: true
      }
    }
    // tile row {
    //   item value {
    //     value: "Renewal Rate"
    //   }
    //   item metric {
    //     value: finance:RevenueRenewalRate * 100
    //     target: 100
    //     view: metric
    //     format: percentage
    //   }
    // }
    tile row {
      item value {
        value: "Growth Rate"
      }
      item metric {
        value: @index.SpendTrend
        target: 100
        view: metriccell
        format: spendtrend
      }
    }
    tile row {
      item value {
        value: "Likelihood To Renew"
      }
      item metric {
        value: average(score(teamcheck:Q2), @daterange.currentPeriodTC)
        view: metriccell
        target: 8
      }
    }
    tile row {
      item value {
        value: "Support Future Needs"
      }
      item metric {
        value: average(score(relationship:Q12), @daterange.currentPeriodRel)
        view: metriccell
        target: 7
      }
    }

  }

  widget keyDrivers #KDAmediumM {

    suppressRule {
      criteria: count(relationship:responseid, (@filter.isPartial OR @filter.isResponded) AND @daterange.currentPeriodRel) = 0
      label: "No responses found"
    }
    label: "Key Drivers"
    size: large
    algorithm: correlation
    importanceLimit: 0.62
    satisfactionLimit: 78
    quadrantTitles: "Improve (High Priority)","Maintain", "Improve (Low Priority)","Watch"
    dependentVariable: relationship:Q1
    independentVariables: relationship:Q4, relationship:Q7, relationship:Q9.1, relationship:Q9.2, relationship:Q9.3, relationship:Q3, relationship:Q12

  }

}

config actionPlanner {
  listPageId: "Initiatives"
  detailsPageId: "InitiativeDetails"
}

page #ConfirmitInitiatives {
  label: "Confirmit Initiatives"

  layoutArea toolbar {
    hide: true
  }
  widget initiativeSummary {
    size: "large"
    items: "totalInitiatives", "myInitiatives", "activeInitiatives", "closedInitiatives"
  }

  widget initiativeList {
    size: "large"
  }

  // widget initiativeProgress {
  //   label: "Initiatives Progress"
  //   size: large
  //   table: apInitiatives:
  //   palette: #82D854,#F0AD4C, #FA5263
  // }

}

page #InitiativeDetails {
  label: "InitiativeDetails"

  hide: true
  widget initiativeDetailSummary {
    size: "large"
  }

  widget initiativeTrend {
    size: "large"
  }

  widget initiativeActions {
    size: "halfwidth"
  }

  widget initiativeNotes {
    size: "halfwidth"
  }
}

page account #Response {
  label: "Response"

  modal: true
  widget contactSurveyResponse {
    view title #defaultSurveyResponseTitle {
    }
    size: medium


    surveyResponseTitle {
      tile title #rt {
        value: contacts:FirstName + " " + contacts:LastName + " - Relationship Survey"
        surveyName: "Relationship Survey"
        view: defaultSurveyResponseTitle
      }
    }

    summary {
      rows: 4
      tile list #list1 {
        item value {
          value: relationship:status
          label: "Status"
        }
        item date {
          value: relationship:interview_start
          label: "Feedback Received"
          format: long
        }
      }
      tile list #list2 {
        item value {
          value: "Relationship Survey"
          label: "Source"
        }
        item value {
          value: relationship:responseid
          label: "Response ID"
        }
      }
    }
 // end of summary

    tab {
      label: "Responses"
      tile list {
        label: " "
        item comment {
          label: "First Name"
          value: contacts:FirstName
        }
        item comment {
          label: "Last Name"
          value: contacts:LastName
        }
        item comment {
          label: "Company name"
          value: SFDCAccounts:Name
        }
        item comment {
          label: "Title"
          value: contacts:Title
        }
        item comment {
          label: "Customer Type"
          value: SFDCAccounts:ClientType
        }
        item comment {
          label: "Role"
          value: contacts:ContactRole
        }
      }
      tile list {
        label: "Key Metrics"
        item bar {
          label: "Likelihood to Recommend"
          value: average(score(relationship:q1))
        }
        item comment {
          label: "Likelihood to Recommend comment"
          value: relationship:Q2
        }
        item bar {
          label: "Satisfaction with Relationship"
          value: average(score(relationship:q4))
        }
        item comment {
          label: "Satisfaction with Relationship comment"
          value: relationship:Q6
        }
        item bar {
          label: "Satisfaction with Technology"
          value: average(score(relationship:q7))
        }
        item comment {
          label: "Satisfaction with Technology comment"
          value: relationship:Q8
        }
      }
      tile list {
        label: "Product"
        item bar {
          label: "Product is reliable"
          value: average(score(relationship:q9.1))
        }
        item bar {
          label: "Product is user friendly"
          value: average(score(relationship:q9.2))
        }
        item bar {
          label: "Product fulfills business needs"
          value: average(score(relationship:q9.3))
        }
      }

      tile list {
        label: "Service"
        item bar {
          label: "Working with Confirmit added value"
          value: average(score(relationship:q3))
        }
        item bar {
          label: "Confirmit can continue to support business needs"
          value: average(score(relationship:q12))
        }
        item comment {
          label: "Why support business needs"
          value: relationship:Q5
        }
        item comment {
          label: "Areas of Improvement"
          value: relationship:Q11
        }
      }
    }
  }
}

//voxpopme
config voxpopme #voxpopmeConfig {
  accountId: 2008
  apiKey: "5df3fb21d0f53ls2rS4o5YFfhZ991GLl "
}

page #TellMeAStory {
  label: "Tell me a story" // - to be added by Tamara on receipt of VoxPopMe login
  widget markdown {
    label: "Tell me a story ... "
    markdown: "[<Ctrl>  &  Click here to record a new video](https://www.confirmit.com/tellmeastory)
   ![picture](https://studio.euro.confirmit.com/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/MRE2EDemo/xzbit.jpg)"

  }

  widget markdown {
    label: "Please note ! "
    markdown: "These videos are confidential. Please do not share any of the videos externally!
    ![picture](https://i.imgflip.com/25nymf.jpg)"

  }


  widget mediaGallery {
    // filter expression {
    //   value: not(feedback:verbatim = "")
    // }
    label: "Videos"
    table: feedback:

    sortBy: feedback:respid
    sortOrder: descending
    size: large
    itemsPerRow: 8
    mediaSource: voxpopmeConfig

    metadata value {
      value: feedback:q8
    }
    metadata value {
      value: feedback:Q1
    }
    metadata value {
      value: feedback:Q2
    }
    metadata value {
      value: feedback:q6
    }
    metadata value {
      value: feedback:q7
    }
    metadata value {
      value: feedback:interview_start
    }
        // voxpopme data
    metadata voxpopme {
      value: "sentimentReadable" // properties from voxpopme REST API response
      label: "Sentiment"
    }
    metadata voxpopme {
      value: "transcripts"
    }
  }
}

page #GiveUsFeedback {
  label: "Give Us Feedback"

  layoutArea toolbar {
    hide: true
  }

  widget markdown {
    size: small
    label: "Your Feedback Is Important. We're listening!"
    markdown: "
[Let Us Know Before You Go](https://survey.euro.confirmit.com/wix/3/p1871616863.aspx)
"
  }

}

page #DrillDown {
  label: "DrillDown"

  modal: true


  widget contactList #hg {
    label: "Response history"
    table: relationship:
    sortColumn: surveyDate
    sortOrder: descending
    size: medium


    view metric #metrics {
      backgroundColorFormatter: backgroundColorFormatter
      valueColorFormatter: valueColorFormatter
      fontSize: small
    }

    column date #inviteDate {
      label: "Request Date"
      value: respondent:smtpstatusDate
      format: dateDefaultFormatter
    }
    column date #surveyDate {
      label: "Response Date"
      value: relationship:interview_start
      format: dateDefaultFormatter
    }

    column value #survey {
      label: "Survey"
      value: "Relationship"
    }

    column metric #ltr {
      label: "LTR"
      value: average(score(relationship:Q1))
      view: metrics
      target: 9
      align: center
    }

    column value #comments {
      label: "Comments"
      value: relationship:Q2
    }

  }
}
