//https://pr.staging.firmglobal.net/apps/editor/201654/page_MainOverview
title "Voice of Guest Dashboard"
//updated: Feb 28, 2024

config hub {
  hub: 12
  numRequests: 4

  dataset survey #surveyDataset {
    publicName: p321993779675 //Delaware North - Master Combined Hub Survey (p321993779675)
    measure filter #filterMeasure_DNListensSurvey {
      value: selected(:survey_pid, @reportConfig.surveypid_dnlistens)
      //value: :survey_name = "DN Listens"
      label: "DN Listens Only"
    }
    measure filter #filterMeasure_ContactRequested {
      value: selected(:CONTACT, "1")
      label: "Contact Req = Yes"
    }
    measure filter #filterMeasure_TeamRecog {
      value: selected(:TEAM_REC, "1")
      label: "Recog = Yes"
    }
    measure filter #filterMeasure_DNListensTravelOnly {
      value: selected(:survey_pid, @reportConfig.surveypid_dnlistens) AND _not(selected(:LocationFinal, @reportConfig.DNListensParkLocations, @reportConfig.DNListensRestaurantLocations))
     // value: :survey_name = "DN Listens" AND _not(IN(:LocationFinal, @reportConfig.DNListensNonTravel))

      label: "DN Listens-Travel locations only"
    }

    measure filter #filterMeasure_DNListensNonTravel {
      value: selected(:survey_pid, @reportConfig.surveypid_dnlistens) AND selected(:LocationFinal, @reportConfig.DNListensNonTravelLocations)
      label: "DN Listens-Non-Travel locations"
    }

    measure filter #filterMeasure_DNListensRestaurants {
      value: selected(:survey_pid, @reportConfig.surveypid_dnlistens) AND selected(:LocationFinal, @reportConfig.DNListensRestaurantLocations)
      label: "DN Listens-Restaurant locations"
    }

    measure filter #filterMeasure_DNListensParks {
      value: selected(:survey_pid, @reportConfig.surveypid_dnlistens) AND selected(:LocationFinal, @reportConfig.DNListensParkLocations)
      label: "DN Listens-Parks locations"
    }

    measure filter #filterMeasure_NPSanswered {
      value: _isnotnull(:NPS) OR _isnotnull(:SAT)
      label: "NPS or OSAT has a value"
    }

    measure filter #filterMeasure_LodgingSurvey {
      value: selected(:survey_pid, @reportConfig.surveypid_lodging)
     // value: :survey_name = "DN Lodging"
      label: "Lodging Only"
    }

    measure filter #filterMeasure_GamingSurvey {
      value: selected(:survey_pid, @reportConfig.surveypid_gaming)
      label: "Gaming Only"
    }


    measure filter #filterMeasure_KSCVCSurvey {
      value: selected(:survey_pid, @reportConfig.surveypid_kscvc)
      label: "Kennedy Space Center"
    }

    measure filter #filterMeasure_ToursSurvey {
      value: selected(:survey_pid, @reportConfig.surveypid_tours)
      label: "Tours Only"
    }

    measure filter #filterMeasure_LizardIslandSurvey {
      value: selected(:survey_pid, @reportConfig.surveypid_lizard)
      label: "Lizard Island Only"
    }

    measure filter #filterMeasure_RatedRestaurant {
      value: _isnotnull(:RESTAURANT_INSERT_TEXT)
      label: "Restaurant Answered"
    }


    measure filter #filterMeasure_Southland_Gaming_Segs {
      value: _isnotnull(:Southland_Gaming_Seg_assign)
      label: "Southland Gaming Segments"
    }

    measure filter #filterMeasure_AustraliaLocations {
      value: selected(:LocationFinal, @reportConfig.AustraliaLocations)
      label: "Australia locations"
    }

    measure filter #filterMeasure_ExcludeAustraliaLocations {
      value: _not(selected(:LocationFinal, @reportConfig.AustraliaLocations))
      label: "Exclude Australia locations"
    }

  }
  dataSet: surveyDataset

//relation needed to connect combined Hub survey with TA survey
//primary key should be combined (i.e. the combined hub survey)
//foreign key should be the TA survey 
  relation oneToOne {
    primaryKey: surveyDataset:survey_rid
    foreignKey: surveyDataset_TA:survey_rid
  }

  //setup for Access Rules
  table accessRules = Studio.DN_Access_Rules
  userProperty claim #UserSegment {// adds a new value on @currentUser object that we can refer to later e.g. in filter
    joinKey: accessRules:UserName// username to match on currently logged in user
    value: accessRules:UserSegment// which corresponding column value we want to use
  }

  userProperty claim #UserLevel {// adds a new value on @currentUser object that we can refer to later e.g. in filter
    joinKey: accessRules:UserName// username to match on currently logged in user
    value: accessRules:UserLevel// which corresponding column value we want to use
  }


  //added for Action Mgmt
  // table amTable = am.CASE
  dataset custom #amTable {
    publicName: am
    defaultTable: CASE
    measure filter #filterMeasure_AMCasesOpen {
      value: selected(amTable:lk_3827, "14869")
      label: "Cases - Open"
    }

    measure filter #filterMeasure_AMCasesInProg {
      value: selected(amTable:lk_3827, "14874")
      label: "Cases - In Progress"
    }
    measure filter #filterMeasure_AMCasesOverdue {
      value: selected(amTable:lk_3827, "14869", "14874") AND amTable:DateDue < GetDate()
      label: "Cases - Overdue"
    }


  }

  variable numeric #daysToClose {
    label: "Days to Close"
    table: amTable:
    value: DiffDay(amTable:DateCreated, IIF(amTable:SystemStatus = "open", GetDate(), amTable:DateClosed))
  }

  variable singleChoice #NPSVal {
    table: surveyDataset:
    value: IIF(score(@reportConfig.nps_qid) >= 9, "A", IIF(score(@reportConfig.nps_qid) >= 7, "B", IIF(score(@reportConfig.nps_qid) >= 0, "C")))
    option code {
      code: "C"
      score: 1
      label: "Detractors"
    }

    option code {
      code: "B"
      score: 2
      label: "Passives"
    }

    option code {
      code: "A"
      score: 3
      label: "Promoters"
    }
  }

  variable singleChoice #RegionRecode {
    table: surveyDataset:
    value: IIF(IN(surveyDataset:REGION, "1"), "US", "Intl")
    option code {
      code: "US"

      label: "U.S."
    }

    option code {
      code: "Intl"

      label: "International"
    }

  }


  dataset custom #Goals_CustomTable {
    publicName: Studio
    defaultTable: DN_Location_Goals
  }
  relation oneToMany {
    primaryKey: Goals_CustomTable:id
    foreignKey: :LocationFinal

  }


   // derived variable/recoding for respondent status
  variable singleChoice #responseStatus {
    table: .respondent:
    label: "Status"
    //value: IIF(survey:status = "Complete", "c", IIF(.respondent:status = "Incomplete", "i", IIF(.respondent:status = "Screened", "s", IIF(.respondent:status = "Quotafull", "q", "n"))))
    value: IIF(.respondent:status = "Complete", "c", IIF(.respondent:status = "Incomplete", "i", IIF(.respondent:smtpStatus = "messageSent", "n", "")))

    option code {
      code: "c"
      label: "Complete"
    }
    option code {
      code: "i"
      label: "Incomplete"
    }
    // option code {
    //   code: "s"
    //   label: "Screened"
    // }
    // option code {
    //   code: "q"
    //   label: "Quota full"
    // }
    option code {
      code: "n"
      label: "Not started"
    }
  } // end variable
  recoding values #sevenPtAgree3cats {

    mapping {
      to: "% Agree (Bottom)"
      from: "'1'..'2'"
    }
    mapping {
      to: "% Agree (Middle)"
      from: "'3'..'5'"
    }
    mapping {
      to: "% Agree (Top)"
      from: "'6'..'7'"
    }
  }

  categorySet #categorySet_meal_rated {
    question: surveyDataset:MEAL_RATED

  }

  // categorySet #categorySet_restaurant_rated {
  //   question: surveyDataset:RESTAURANT_INSERT

  // }

  categorySet #categorySet_premium_exp_rated {
    question: surveyDataset:PREMIUM_INSERT

  }


  categorySet #categorySet_shop_rated {
    question: surveyDataset:SHOPS_INSERT

  }

  categorySet #categorySet_attraction_rated {
    question: surveyDataset:ATTRACT_INSERT

  }

  //define reusable selector lists
  valueSet #valueSet_date_ranges_1 {
		// item {
		// 	label: "Daily"

		// 	value:  {
		// 		selectBreakdownBy: "calendarDate"
		// 		selectFilter: InDay(@reportConfig.intvdate, -30, 0)
		// 	}
		// }
		// item {
		// 	label: "Weekly"

		// 	value:  {
		// 		selectBreakdownBy: "calendarWeek"
		// 		selectFilter: InDay(@reportConfig.intvdate, -84, 0) //84 days is 12 weeks
		// 	}
		// }
    item {
      label: "Monthly"

      value:  {
        selectBreakdownBy: "calendarMonth"
        selectFilter: InMonth(@reportConfig.intvdate, -11, 0)
        selectStart: "-12 month"
      }
    }
    item {
      label: "Quarterly"

      value:  {
        selectBreakdownBy: "calendarQuarter"
        selectFilter: InQuarter(@reportConfig.intvdate, -7, 0)
        selectStart: "-7 quarter"
      }
    }
    item {
      label: "Yearly"

      value:  {
        selectBreakdownBy: "Year"
        selectFilter: InYear(@reportConfig.intvdate, -2, 0)
        selectStart: "-2 year"
      }
    }

  } // end valueSet
  valueSet #valueSet_date_ranges_RR {
    // item {
    //   label: "Daily"

    //   value:  {
    //     selectBreakdownBy: "calendarDate"
    //     selectFilter: InDay(@reportConfig.InvitedDate, -14, 0)
    //   }
    // }
    // item {
    //   label: "Weekly"

    //   value:  {
    //     selectBreakdownBy: "calendarWeek"
    //     selectFilter: InDay(@reportConfig.InvitedDate, -42, 0) //42 days is 6 weeks, 84 days is 12 weeks
    //   }
    // }
    item {
      label: "Monthly"

      value:  {
        selectBreakdownBy: "calendarMonth"
        selectFilter: InMonth(@reportConfig.InvitedDate, -11, 0)

      }
    }
    item {
      label: "Quarterly"

      value:  {
        selectBreakdownBy: "calendarQuarter"
        selectFilter: InQuarter(@reportConfig.InvitedDate, -7, 0)

      }
    }
    item {
      label: "Yearly"

      value:  {
        selectBreakdownBy: "Year"
        selectFilter: InYear(@reportConfig.InvitedDate, -2, 0)

      }
    }

  } // end valueSet
  valueSet #valueSet_lodging_locations {

    item {
      label: "Lodging locations"
      value: "Lodging"
    }

    item {
      label: "The Lodge at Tenaya"
      value: "474A"
    }

    item {
      label: "The Cottages at Tenaya"
      value: "474B"
    }

    item {
      label: "The Explorer Cabins at Tenaya"
      value: "474C"
    }

    item {
      label: "Yavapai Lodge - Grand Canyon National Park"
      value: "63108"
    }

    item {
      label: "Trailer Village RV Park - Grand Canyon National Park"
      value: "63275"
    }

    item {
      label: "Skyland Resort - Shenandoah National Park"
      value: "58867"
    }

    item {
      label: "Big Meadows Lodge - Shenandoah National Park"
      value: "58866"
    }

    // item {
    //   label: "Lewis Mountain Cabins - Shenandoah National Park"
    //   value: "58865"
    // }

    item {
      label: "The Lodge at Geneva on the Lake"
      value: "22005A"
    }

    item {
      label: "The Cottages at Geneva on the Lake"
      value: "22005B"
    }

    // item {
    //   label: "Cedar Grove Lodge - Kings Canyon National Park"
    //   value: "59988"
    // }

    item {
      label: "Grant Grove Cabins - Kings Canyon National Park"
      value: "59989B"
    }

    item {
      label: "John Muir Lodge - Kings Canyon National Park"
      value: "59989A"
    }

    item {
      label: "Wuksachi Lodge - Sequoia National Park"
      value: "404"
    }

    item {
      label: "Kalaloch Lodge"
      value: "58148"
    }

    item {
      label: "The Explorer Cabins - Yellowstone"
      value: "59396"
    }

    item {
      label: "Gray Wolf Inn & Suites - Yellowstone"
      value: "28577"
    }

    item {
      label: "Yellowstone Park Hotel"
      value: "28578"
    }

    item {
      label: "Peaks of Otter"
      value: "59841"
    }

    item {
      label: "The Gideon Putnam"
      value: "139"
    }

  } // end valueSet valueSet_lodging_locations
  valueSet #valueSet_gaming_locations {

    item {
      label: "Gaming locations"
      value:  {
        selectCode: "Gaming"
        selectHotelCode: ""
        selectFilter: true
      }
    }

    // item {
    //   label: "Catawba Two Kings Casino"
    //   value: "TK"
    // }

    // item {
    //   label: "Daytona Beach Racing and Card Club"
    //   value: "DB"
    // }	

    item {
      label: "Finger Lakes Gaming"
      value:  {
        selectCode: "FL"
        selectHotelCode: ""
        selectFilter: selected(:LocationFinal, "FL")
      }
    }

    item {
      label: "Gate City Casino"
      value:  {
        selectCode: "BB"
        selectHotelCode: ""
        selectFilter: selected(:LocationFinal, "BB")
      }
    }

    item {
      label: "Hamburg Gaming"
      value:  {
        selectCode: "HB"
        selectHotelCode: ""
        selectFilter: selected(:LocationFinal, "HB")
      }
    }

    item {
      label: "Mardi Gras Casino & Resort"
      value:  {
        selectCode: "MG"
        selectHotelCode: "7689"
        selectFilter: selected(:LocationFinal, "MG", "7689")

      }

    }

    // item {
    //   label: "Mardi Gras Casino & Resort Hotel"
    //   value: "7689"
    // }

    item {
      label: "Miami Valley Gaming"
      value:  {
        selectCode: "MVG"
        selectHotelCode: ""
        selectFilter: selected(:LocationFinal, "MVG")
      }
    }

    // item {
    //   label: "Mindil Beach Casino Resort"
    //   value: "MBCR"
    // }

    // item {
    //   label: "Mindil Beach Casino Resort Hotel"
    //   value: "40765"
    // }

    // item {
    //   label: "Orange City Racing and Card Club"
    //   value: "OC"
    // }	

    item {
      label: "Southland Casino Resort"
      value:  {
        selectCode: "SL"
        selectHotelCode: "38344"
        selectFilter: selected(:LocationFinal, "MG", "38344")

      }
    }

    // item {
    //   label: "Southland Casino Hotel"
    //   value: "38344"
    // }

    item {
      label: "Wheeling Island Casino Resort"
      value:  {
        selectCode: "WI"
        selectHotelCode: "51559"
        selectFilter: selected(:LocationFinal, "WI", "51559")

      }
    }

    // item {
    //   label: "Wheeling Island Hotel - Casino - Racetrack"
    //   value: "51559"
    // }

  } // end valueSet valueSet_gaming_locations
  valueSet #valueSet_tours_locations {

    item {
      label: "Tours locations"
      value: "Tours"
    }

    item {
      label: "Nova Guides at Camp Hale"
      value: "Nova_Guides_1"
    }

    item {
      label: "Shenandoah National Park Tours"
      value: "Shenandoah_Tours_1"
    }

    item {
      label: "Yellowstone Vacation Tours - West Yellowstone"
      value: "Yellowstone_Tours_1"
    }

    item {
      label: "Yosemite 360 Tours"
      value: "Yosemite_Tours_1"
    }

  }

  valueSet #valueSet_australia_locations {

    item {
      label: "Australia locations"
      value: "Australia"
    }

    item {
      label: "Lizard Island"
      value: "51906"
    }
  }

  valueSet #valueSet_date_ranges {

		// item {
		// 	label: "Daily"

		// 	value:  {
		// 		selectBreakdownBy: "calendarDate"
		// 		selectFilter: InDay(@reportConfig.intvdate, -30, 0)
		// 	}
		// }
		// item {
		// 	label: "Weekly"

		// 	value:  {
		// 		selectBreakdownBy: "calendarWeek"
		// 		selectFilter: InDay(@reportConfig.intvdate, -84, 0) //84 days is 12 weeks
		// 	}
		// }
    item {
      label: "Monthly"

      value:  {
        selectBreakdownBy: "calendarMonth"
        selectFilter: InMonth(@reportConfig.intvdate_ta, -11, 0)
      }
    }
    item {
      label: "Quarterly"

      value:  {
        selectBreakdownBy: "calendarQuarter"
        selectFilter: InQuarter(@reportConfig.intvdate_ta, -19, 0)

      }
    }
    item {
      label: "Yearly"

      value:  {
        selectBreakdownBy: "Year"
        selectFilter: InYear(@reportConfig.intvdate_ta, -4, 0)

      }
    }

  } // end valueSet	
  valueSet #valueSet_hierarchy_views {
    item {
      label: "Hierarchical View"
      value: 1
    }
    item {
      label: "Flat View"
      value: 2
    }
  } // end valueSet	 
  reportingHierarchy selfRefLookup #SitesHierarchy {
    source: :LocationFinal
    label: "Delaware North - Main Hierarchy"
  }
  reportingHierarchy selfRefLookup #SitesHierarchySimplified {
    source: :LocationSimplified
    label: "Delaware North - Simplified Hierarchy"
    showBreadcrumb: true
  }

  reportingHierarchy surveyBased #LocationsBySurveyHierarchy {
    label: "Locations By Survey"
    level #level1 {
      value: surveyDataset.respondent:survey_pid

    }
    level #level2 {
      value: surveyDataset.respondent:LocationName

    }
  }
  reportingHierarchy surveyBased #RestaurantHierarchy {
    level #level1 {
      value: surveyDataset:LocationName
    }
    label: "Restaurant Hierarchy"
    level #level2 {
      value: surveyDataset:RESTAURANT_INSERT_TEXT
    }
  }

  //begin TA dataset
  dataset survey #surveyDataset_TA {
    publicName: p438345471506
    variable singleChoice #NPSVal {
      table: surveyDataset_TA:
      value: IIF(score(@reportConfig.nps_qid_ta) >= 9, "A", IIF(score(@reportConfig.nps_qid_ta) >= 7, "B", IIF(score(@reportConfig.nps_qid_ta) >= 0, "C")))
      option code {
        code: "C"
        score: 1
        label: "Detractors"
      }

      option code {
        code: "B"
        score: 2
        label: "Passives"
      }

      option code {
        code: "A"
        score: 3
        label: "Promoters"
      }
    }
  }
  dataset textAnalytics #textAnalyticsDataset_Lodging {
    publicName: TextAnalytics_p438345471506_4072
    table responses = p438345471506.response:
    propagateFilter #propagateFilter_1 {
      from: .model:
      to: .categoryScore:
    }
    propagateFilter #propagateFilter_2 {
      from: .categoryScore:
      to: .overallScore:
    }
    propagateFilter #propagateFilter_3 {
      from: .overallScore:
      to: .responses:
    }
    propagateFilter #propagateFilter_4 {
      from: .overallScore:
      to: .analysisRecord:
    }
    variable singleChoice #PosNegNeutralGroupsOverallSentiment {
      table: textAnalyticsDataset_Lodging.overallScore:
      value: iif(textAnalyticsDataset_Lodging.overallScore:score > 0, "positive", iif(textAnalyticsDataset_Lodging.overallScore:score = 0, "neutral", iif(textAnalyticsDataset_Lodging.overallScore:score < 0, "negative")))

      option code {
        code: "positive"
        label: "Positive"
        score: 3
      }

      option code {
        code: "neutral"
        label: "Neutral"
        score: 2
      }

      option code {
        code: "negative"
        label: "Negative"
        score: 1
      }

    }

    variable singleChoice #PosNegNeutralGroups {
      table: textAnalyticsDataset_Lodging.categoryScore:
      value: iif(textAnalyticsDataset_Lodging.categoryScore:score > 0, "positive", iif(textAnalyticsDataset_Lodging.categoryScore:score = 0, "neutral", iif(textAnalyticsDataset_Lodging.categoryScore:score < 0, "negative")))

      option code {
        code: "positive"
        label: "Positive"
        score: 3
      }

      option code {
        code: "neutral"
        label: "Neutral"
        score: 2
      }

      option code {
        code: "negative"
        label: "Negative"
        score: 1
      }

    }

    reportingHierarchy selfRefCustom #categoryHierarchy_Lodging {
      label: "Categories model"
      mode: "direct"
      parent: textAnalyticsDataset_Lodging.model:parent
      nodeLabel: textAnalyticsDataset_Lodging.model:label
    }

 //Overall measures
// overallCount() - Number of overall sentiments
// overallAverage() - Average overall sentiment
// overallResponseBase() - Number of responses in overall sentiments
// overallRespondentBasePercent() - Percentage of respondents in overall sentiments
// overallCommentsBase() - Number of comments with overall sentiments
// overallCommentsPercent() - Percentage of comments with overall sentiments
// overallPositiveCount() - Count of positive overall sentiments
// overallPositivePercent() - Percentage of positive overall sentiments
// overallNeutralCount() - Count of neutral overall sentiment
// overallNeutralPercent() - Percentage of neutral overall sentiments
// overallNegativeCount() - Count of negative overall sentiments
// overallNegativePercent() - Percentage of negative overall sentiments

//Categories measures
// categoryCount() - Number of categories
// categoryAverage() - Average category sentiment
// categoryResponseBase() - Number of responses within category
// categoryRespondentBasePercent() - Percentage of respondents within category
// categoryCommentsBase() - Number of comments categorised
// categoryCommentsPercent() - Percentage of comments categorised
// categoryPositiveCount() - Count of positive category sentiments
// categoryPositivePercent() - Percentage of positive category sentiments
// categoryNeutralCount() - Count of neutral category sentiments
// categoryNeutralPercent() - Percentage of neutral category sentiments
// categoryNegativeCount() - Count of negative category sentiments
// categoryNegativePercent() - Percentage of negative category sentiments


    //CATEGORY LEVEL
    measure custom #categoryCountTASet1 { //default measure here just in case
      value: count(textAnalyticsDataset_Lodging.categoryScore:)
      label: "Number of comments by category"
    }
    measure custom #categoryAverageTASet1 { //default measure here just in case
      value: average(textAnalyticsDataset_Lodging.categoryScore:score)
      label: "Average category sentiment"
    }
    measure custom #categoryResponseBaseTASet1 { //default measure here just in case
      value: countDistinct(textAnalyticsDataset_Lodging.categoryScore:responseId)
      label: "Number of responses within category"
    }
    measure custom #respondentsAllCategoriesPositiveCountTASet1 {
      label: "Number of respondents that are positive through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Lodging.responses:), textAnalyticsDataset_Lodging.categoryScore:), avg(textAnalyticsDataset_Lodging.categoryScore:score, true, textAnalyticsDataset_Lodging.responses:) > 0.25)
    }
    measure custom #respondentsAllCategoriesNeutralCountTASet1 {
      label: "Number of respondents that are neutral through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Lodging.responses:), textAnalyticsDataset_Lodging.categoryScore:), avg(textAnalyticsDataset_Lodging.categoryScore:score, true, textAnalyticsDataset_Lodging.responses:) = 0)
    }
    measure custom #respondentsAllCategoriesNegativeCountTASet1 {
      label: "Number of respondents that are negative through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Lodging.responses:), textAnalyticsDataset_Lodging.categoryScore:), avg(textAnalyticsDataset_Lodging.categoryScore:score, true, textAnalyticsDataset_Lodging.responses:) < -0.25)
    }

    //COMMENT LEVEL

    measure custom #commentsOverallCountTASet1 {
      label: "Number of comments overall"
      value: count(textAnalyticsDataset_Lodging.overallScore:responseid)
    }
    measure custom #commentsOverallPositiveCountTASet1 {
      label: "Number of positive comments overall"
      value: count(textAnalyticsDataset_Lodging.overallScore:responseid, textAnalyticsDataset_Lodging.overallScore:score > 0)
    }

    measure custom #commentsOverallNeutralCountTASet1 {
      label: "Number of neutral comments overall"
      value: count(textAnalyticsDataset_Lodging.overallScore:responseid, textAnalyticsDataset_Lodging.overallScore:score = 0)
    }

    measure custom #commentsOverallNegativeCountTASet1 {
      label: "Number of negative comments overall"
      value: count(textAnalyticsDataset_Lodging.overallScore:responseid, textAnalyticsDataset_Lodging.overallScore:score < 0)
    }

    measure custom #respondentsOverallPositiveCountTASet1 {
      label: "Number of respondents that are overall positive"
      value: countIf(average(textAnalyticsDataset_Lodging.overallScore:score, true, textAnalyticsDataset_Lodging.responses:) > 0)
    }
    measure custom #respondentsOverallNeutralCountTASet1 {
      label: "Number of respondents that are overall neutral"
      value: countIf(average(textAnalyticsDataset_Lodging.overallScore:score, true, textAnalyticsDataset_Lodging.responses:) = 0)
    }
    measure custom #respondentsOverallNegativeCountTASet1 {
      label: "Number of respondents that are overall negative"
      value: countIf(average(textAnalyticsDataset_Lodging.overallScore:score, true, textAnalyticsDataset_Lodging.responses:) < 0)
    }

    //OVERALL LEVEL
    measure custom #overallAverageTASet1 { //default measure here just in case
      value: average(textAnalyticsDataset_Lodging.overallScore:score)
      label: "Average overall sentiment"
    }
    measure custom #overallResponseBaseTASet1 { //default measure here just in case
      value: countDistinct(textAnalyticsDataset_Lodging.overallScore:responseId)
      label: "Number of respondents in overall sentiments"
    }
    measure custom #overallPositiveAverageTASet1 {
      label: "Average positive overall sentiment"
      value: avg(textAnalyticsDataset_Lodging.overallScore:score, textAnalyticsDataset_Lodging.overallScore:score > 0)
    }
    measure custom #overallNegativeAverageTASet1 {
      label: "Average negative overall sentiment"
      value: avg(textAnalyticsDataset_Lodging.overallScore:score, textAnalyticsDataset_Lodging.overallScore:score < 0)
    }
    measure custom #overallPositivePercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Lodging.overallScore:overallSentimentGroup, "positive")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #overallNeutralPercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Lodging.overallScore:overallSentimentGroup, "neutral")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #overallNegativePercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Lodging.overallScore:overallSentimentGroup, "negative")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #percentageOfCommentsTASet1 {
      label: "Percentage of overall distinct comments"
      value: 100 * countDistinct(demote(recordId(textAnalyticsDataset_Lodging.overallScore:), textAnalyticsDataset_Lodging.categoryScore:)) / count(textAnalyticsDataset_Lodging.overallScore:, true, "__top")
    }

  } // end textAnalyticsDataset_Lodging
  dataset textAnalytics #textAnalyticsDataset_Gaming {
    publicName: TextAnalytics_p438345471506_4089
    table responses = p438345471506.response:
    propagateFilter #propagateFilter_1 {
      from: .model:
      to: .categoryScore:
    }
    propagateFilter #propagateFilter_2 {
      from: .categoryScore:
      to: .overallScore:
    }
    propagateFilter #propagateFilter_3 {
      from: .overallScore:
      to: .responses:
    }
    propagateFilter #propagateFilter_4 {
      from: .overallScore:
      to: .analysisRecord:
    }
    variable singleChoice #PosNegNeutralGroupsOverallSentiment {
      table: textAnalyticsDataset_Gaming.overallScore:
      value: iif(textAnalyticsDataset_Gaming.overallScore:score > 0, "positive", iif(textAnalyticsDataset_Gaming.overallScore:score = 0, "neutral", iif(textAnalyticsDataset_Gaming.overallScore:score < 0, "negative")))

      option code {
        code: "positive"
        label: "Positive"
        score: 3
      }

      option code {
        code: "neutral"
        label: "Neutral"
        score: 2
      }

      option code {
        code: "negative"
        label: "Negative"
        score: 1
      }

    }

    variable singleChoice #PosNegNeutralGroups {
      table: textAnalyticsDataset_Gaming.categoryScore:
      value: iif(textAnalyticsDataset_Gaming.categoryScore:score > 0, "positive", iif(textAnalyticsDataset_Gaming.categoryScore:score = 0, "neutral", iif(textAnalyticsDataset_Gaming.categoryScore:score < 0, "negative")))

      option code {
        code: "positive"
        label: "Positive"
        score: 3
      }

      option code {
        code: "neutral"
        label: "Neutral"
        score: 2
      }

      option code {
        code: "negative"
        label: "Negative"
        score: 1
      }

    }

    reportingHierarchy selfRefCustom #categoryHierarchy_Gaming {
      label: "Categories model"
      mode: "direct"
      parent: textAnalyticsDataset_Gaming.model:parent
      nodeLabel: textAnalyticsDataset_Gaming.model:label
    }

 //Overall measures
// overallCount() - Number of overall sentiments
// overallAverage() - Average overall sentiment
// overallResponseBase() - Number of responses in overall sentiments
// overallRespondentBasePercent() - Percentage of respondents in overall sentiments
// overallCommentsBase() - Number of comments with overall sentiments
// overallCommentsPercent() - Percentage of comments with overall sentiments
// overallPositiveCount() - Count of positive overall sentiments
// overallPositivePercent() - Percentage of positive overall sentiments
// overallNeutralCount() - Count of neutral overall sentiment
// overallNeutralPercent() - Percentage of neutral overall sentiments
// overallNegativeCount() - Count of negative overall sentiments
// overallNegativePercent() - Percentage of negative overall sentiments

//Categories measures
// categoryCount() - Number of categories
// categoryAverage() - Average category sentiment
// categoryResponseBase() - Number of responses within category
// categoryRespondentBasePercent() - Percentage of respondents within category
// categoryCommentsBase() - Number of comments categorised
// categoryCommentsPercent() - Percentage of comments categorised
// categoryPositiveCount() - Count of positive category sentiments
// categoryPositivePercent() - Percentage of positive category sentiments
// categoryNeutralCount() - Count of neutral category sentiments
// categoryNeutralPercent() - Percentage of neutral category sentiments
// categoryNegativeCount() - Count of negative category sentiments
// categoryNegativePercent() - Percentage of negative category sentiments


    //CATEGORY LEVEL
    measure custom #categoryCountTASet1 { //default measure here just in case
      value: count(textAnalyticsDataset_Gaming.categoryScore:)
      label: "Number of comments by category"
    }
    measure custom #categoryAverageTASet1 { //default measure here just in case
      value: average(textAnalyticsDataset_Gaming.categoryScore:score)
      label: "Average category sentiment"
    }
    measure custom #categoryResponseBaseTASet1 { //default measure here just in case
      value: countDistinct(textAnalyticsDataset_Gaming.categoryScore:responseId)
      label: "Number of responses within category"
    }
    measure custom #respondentsAllCategoriesPositiveCountTASet1 {
      label: "Number of respondents that are positive through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Gaming.responses:), textAnalyticsDataset_Gaming.categoryScore:), avg(textAnalyticsDataset_Gaming.categoryScore:score, true, textAnalyticsDataset_Gaming.responses:) > 0.25)
    }
    measure custom #respondentsAllCategoriesNeutralCountTASet1 {
      label: "Number of respondents that are neutral through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Gaming.responses:), textAnalyticsDataset_Gaming.categoryScore:), avg(textAnalyticsDataset_Gaming.categoryScore:score, true, textAnalyticsDataset_Gaming.responses:) = 0)
    }
    measure custom #respondentsAllCategoriesNegativeCountTASet1 {
      label: "Number of respondents that are negative through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Gaming.responses:), textAnalyticsDataset_Gaming.categoryScore:), avg(textAnalyticsDataset_Gaming.categoryScore:score, true, textAnalyticsDataset_Gaming.responses:) < -0.25)
    }

    //COMMENT LEVEL

    measure custom #commentsOverallCountTASet1 {
      label: "Number of comments overall"
      value: count(textAnalyticsDataset_Gaming.overallScore:responseid)
    }
    measure custom #commentsOverallPositiveCountTASet1 {
      label: "Number of positive comments overall"
      value: count(textAnalyticsDataset_Gaming.overallScore:responseid, textAnalyticsDataset_Gaming.overallScore:score > 0)
    }

    measure custom #commentsOverallNeutralCountTASet1 {
      label: "Number of neutral comments overall"
      value: count(textAnalyticsDataset_Gaming.overallScore:responseid, textAnalyticsDataset_Gaming.overallScore:score = 0)
    }

    measure custom #commentsOverallNegativeCountTASet1 {
      label: "Number of negative comments overall"
      value: count(textAnalyticsDataset_Gaming.overallScore:responseid, textAnalyticsDataset_Gaming.overallScore:score < 0)
    }

    measure custom #respondentsOverallPositiveCountTASet1 {
      label: "Number of respondents that are overall positive"
      value: countIf(average(textAnalyticsDataset_Gaming.overallScore:score, true, textAnalyticsDataset_Gaming.responses:) > 0)
    }
    measure custom #respondentsOverallNeutralCountTASet1 {
      label: "Number of respondents that are overall neutral"
      value: countIf(average(textAnalyticsDataset_Gaming.overallScore:score, true, textAnalyticsDataset_Gaming.responses:) = 0)
    }
    measure custom #respondentsOverallNegativeCountTASet1 {
      label: "Number of respondents that are overall negative"
      value: countIf(average(textAnalyticsDataset_Gaming.overallScore:score, true, textAnalyticsDataset_Gaming.responses:) < 0)
    }

    //OVERALL LEVEL
    measure custom #overallAverageTASet1 { //default measure here just in case
      value: average(textAnalyticsDataset_Gaming.overallScore:score)
      label: "Average overall sentiment"
    }
    measure custom #overallResponseBaseTASet1 { //default measure here just in case
      value: countDistinct(textAnalyticsDataset_Gaming.overallScore:responseId)
      label: "Number of respondents in overall sentiments"
    }
    measure custom #overallPositiveAverageTASet1 {
      label: "Average positive overall sentiment"
      value: avg(textAnalyticsDataset_Gaming.overallScore:score, textAnalyticsDataset_Gaming.overallScore:score > 0)
    }
    measure custom #overallNegativeAverageTASet1 {
      label: "Average negative overall sentiment"
      value: avg(textAnalyticsDataset_Gaming.overallScore:score, textAnalyticsDataset_Gaming.overallScore:score < 0)
    }
    measure custom #overallPositivePercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Gaming.overallScore:overallSentimentGroup, "positive")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #overallNeutralPercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Gaming.overallScore:overallSentimentGroup, "neutral")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #overallNegativePercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Gaming.overallScore:overallSentimentGroup, "negative")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #percentageOfCommentsTASet1 {
      label: "Percentage of overall distinct comments"
      value: 100 * countDistinct(demote(recordId(textAnalyticsDataset_Gaming.overallScore:), textAnalyticsDataset_Gaming.categoryScore:)) / count(textAnalyticsDataset_Gaming.overallScore:, true, "__top")
    }

  } // end textAnalyticsDataset_Gaming
  dataset textAnalytics #textAnalyticsDataset_Dining {
    publicName: TextAnalytics_p438345471506_3561
    table responses = p438345471506.response:
    propagateFilter #propagateFilter {
      from: .model:
      to: .categoryScore:
    }
    propagateFilter #propagateFilter_2 {
      from: .categoryScore:
      to: .overallScore:
    }
    propagateFilter #propagateFilter_3 {
      from: .overallScore:
      to: .responses:
    }
    propagateFilter {
      from: .overallScore:
      to: .analysisRecord:
    }

    reportingHierarchy selfRefCustom #categoryHierarchy_Dining {
      label: "Categories model"
      mode: "direct"
      parent: textAnalyticsDataset_Dining.model:parent
      nodeLabel: textAnalyticsDataset_Dining.model:label
    }



    variable singleChoice #PosNegNeutralGroupsOverallSentiment {
      table: textAnalyticsDataset_Dining.overallScore:
      value: iif(textAnalyticsDataset_Dining.overallScore:score > 0, "positive", iif(textAnalyticsDataset_Dining.overallScore:score = 0, "neutral", iif(textAnalyticsDataset_Dining.overallScore:score < 0, "negative")))

      option code {
        code: "positive"
        label: "Positive"
        score: 3
      }

      option code {
        code: "neutral"
        label: "Neutral"
        score: 2
      }

      option code {
        code: "negative"
        label: "Negative"
        score: 1
      }

    }

    variable singleChoice #PosNegNeutralGroups {
      table: textAnalyticsDataset_Dining.categoryScore:
      value: iif(textAnalyticsDataset_Dining.categoryScore:score > 0, "positive", iif(textAnalyticsDataset_Dining.categoryScore:score = 0, "neutral", iif(textAnalyticsDataset_Dining.categoryScore:score < 0, "negative")))

      option code {
        code: "positive"
        label: "Positive"
        score: 3
      }

      option code {
        code: "neutral"
        label: "Neutral"
        score: 2
      }

      option code {
        code: "negative"
        label: "Negative"
        score: 1
      }

    }

//Overall measures
// overallCount() - Number of overall sentiments
// overallAverage() - Average overall sentiment
// overallResponseBase() - Number of responses in overall sentiments
// overallRespondentBasePercent() - Percentage of respondents in overall sentiments
// overallCommentsBase() - Number of comments with overall sentiments
// overallCommentsPercent() - Percentage of comments with overall sentiments
// overallPositiveCount() - Count of positive overall sentiments
// overallPositivePercent() - Percentage of positive overall sentiments
// overallNeutralCount() - Count of neutral overall sentiment
// overallNeutralPercent() - Percentage of neutral overall sentiments
// overallNegativeCount() - Count of negative overall sentiments
// overallNegativePercent() - Percentage of negative overall sentiments

//Categories measures
// categoryCount() - Number of categories
// categoryAverage() - Average category sentiment
// categoryResponseBase() - Number of responses within category
// categoryRespondentBasePercent() - Percentage of respondents within category
// categoryCommentsBase() - Number of comments categorised
// categoryCommentsPercent() - Percentage of comments categorised
// categoryPositiveCount() - Count of positive category sentiments
// categoryPositivePercent() - Percentage of positive category sentiments
// categoryNeutralCount() - Count of neutral category sentiments
// categoryNeutralPercent() - Percentage of neutral category sentiments
// categoryNegativeCount() - Count of negative category sentiments
// categoryNegativePercent() - Percentage of negative category sentiments


    //CATEGORY LEVEL
    measure custom #categoryCountTASet1 { //default measure here just in case
      value: count(textAnalyticsDataset_Dining.categoryScore:)
      label: "Number of comments by category"
    }
    measure custom #categoryAverageTASet1 { //default measure here just in case
      value: average(textAnalyticsDataset_Dining.categoryScore:score)
      label: "Average category sentiment"
    }
    measure custom #categoryResponseBaseTASet1 { //default measure here just in case
      value: countDistinct(textAnalyticsDataset_Dining.categoryScore:responseId)
      label: "Number of responses within category"
    }
    measure custom #respondentsAllCategoriesPositiveCountTASet1 {
      label: "Number of respondents that are positive through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Dining.responses:), textAnalyticsDataset_Dining.categoryScore:), avg(textAnalyticsDataset_Dining.categoryScore:score, true, textAnalyticsDataset_Dining.responses:) > 0.25)
    }
    measure custom #respondentsAllCategoriesNeutralCountTASet1 {
      label: "Number of respondents that are neutral through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Dining.responses:), textAnalyticsDataset_Dining.categoryScore:), avg(textAnalyticsDataset_Dining.categoryScore:score, true, textAnalyticsDataset_Dining.responses:) = 0)
    }
    measure custom #respondentsAllCategoriesNegativeCountTASet1 {
      label: "Number of respondents that are negative through ALL categories"
      value: countDistinct(demote(recordId(textAnalyticsDataset_Dining.responses:), textAnalyticsDataset_Dining.categoryScore:), avg(textAnalyticsDataset_Dining.categoryScore:score, true, textAnalyticsDataset_Dining.responses:) < -0.25)
    }

    //COMMENT LEVEL

    measure custom #commentsOverallCountTASet1 {
      label: "Number of comments overall"
      value: count(textAnalyticsDataset_Dining.overallScore:responseid)
    }
    measure custom #commentsOverallPositiveCountTASet1 {
      label: "Number of positive comments overall"
      value: count(textAnalyticsDataset_Dining.overallScore:responseid, textAnalyticsDataset_Dining.overallScore:score > 0)
    }

    measure custom #commentsOverallNeutralCountTASet1 {
      label: "Number of neutral comments overall"
      value: count(textAnalyticsDataset_Dining.overallScore:responseid, textAnalyticsDataset_Dining.overallScore:score = 0)
    }

    measure custom #commentsOverallNegativeCountTASet1 {
      label: "Number of negative comments overall"
      value: count(textAnalyticsDataset_Dining.overallScore:responseid, textAnalyticsDataset_Dining.overallScore:score < 0)
    }

    measure custom #respondentsOverallPositiveCountTASet1 {
      label: "Number of respondents that are overall positive"
      value: countIf(average(textAnalyticsDataset_Dining.overallScore:score, true, textAnalyticsDataset_Dining.responses:) > 0)
    }
    measure custom #respondentsOverallNeutralCountTASet1 {
      label: "Number of respondents that are overall neutral"
      value: countIf(average(textAnalyticsDataset_Dining.overallScore:score, true, textAnalyticsDataset_Dining.responses:) = 0)
    }
    measure custom #respondentsOverallNegativeCountTASet1 {
      label: "Number of respondents that are overall negative"
      value: countIf(average(textAnalyticsDataset_Dining.overallScore:score, true, textAnalyticsDataset_Dining.responses:) < 0)
    }

    //OVERALL LEVEL
    measure custom #overallAverageTASet1 { //default measure here just in case
      value: average(textAnalyticsDataset_Dining.overallScore:score)
      label: "Average overall sentiment"
    }
    measure custom #overallResponseBaseTASet1 { //default measure here just in case
      value: countDistinct(textAnalyticsDataset_Dining.overallScore:responseId)
      label: "Number of respondents in overall sentiments"
    }
    measure custom #overallPositiveAverageTASet1 {
      label: "Average positive overall sentiment"
      value: avg(textAnalyticsDataset_Dining.overallScore:score, textAnalyticsDataset_Dining.overallScore:score > 0)
    }
    measure custom #overallNegativeAverageTASet1 {
      label: "Average negative overall sentiment"
      value: avg(textAnalyticsDataset_Dining.overallScore:score, textAnalyticsDataset_Dining.overallScore:score < 0)
    }
    measure custom #overallPositivePercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Dining.overallScore:overallSentimentGroup, "positive")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #overallNeutralPercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Dining.overallScore:overallSentimentGroup, "neutral")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #overallNegativePercentTASet1 { //default measure here just in case
      value: PercentageOfAnswers(textAnalyticsDataset_Dining.overallScore:overallSentimentGroup, "negative")
      label: "Percentage of positive overall sentiments"
    }
    measure custom #percentageOfCommentsTASet1 {
      label: "Percentage of overall distinct comments"
      value: 100 * countDistinct(demote(recordId(textAnalyticsDataset_Dining.overallScore:), textAnalyticsDataset_Dining.categoryScore:)) / count(textAnalyticsDataset_Dining.overallScore:, true, "__top")
    }

//measure filters for TA



  } // end textAnalyticsDataset_Dining
  dataset cases #cases {
    publicName: am
  }
} // end config hub
reportBase #reportBase {
  rule nodesHM #nodesHMRule {
    reportingHierarchy: SitesHierarchy
    //mode: permission
    mode: permission
  }
  rule reportingPeriod #reportingPeriodRule {
    defaultPeriod: "0 year"

  }
}

config queryOptions {
  // added automatically during report creation
  boolNullsAsFalse: false
  explicitLevelAggregation: true


  optimization {
    UseHashJoinHint: "true"
  //  useCrossApplyUnpivot: "true"
  }

}

config layout #layoutConfig {
  horizontalAlignmentMode: "fourColumnsCentered"
}

layoutArea toolbar {
  useDynamicFilters: true
  // filter reportingHierarchy #reportingHierarchyFilter {
  //   reportingHierarchy: SitesHierarchy
  // }
  filter reportingPeriod #reportingPeriodFilter {
    label: "Reporting Period"
  }
  // filter reportingHierarchy #f_SitesHierarchy {
  //   reportingHierarchy: SitesHierarchy
  //   label: "Locations"
  // }

  filter multiselect #f_Location {
    optionsFrom: surveyDataset:LocationName
    label: "Location"

  }

  filter multiselect #f_Surveys {
    optionsFrom: surveyDataset:survey_name
    label: "Survey Name"
  }

  filter multiselect #f_NPS {
    optionsFrom: surveyDataset:NPSVal
    label: "NPS Groups"
  }

  filter multiselect #f_DNListens_SurveyType {
    optionsFrom: surveyDataset:SurveyType
    label: "Survey Type (DN Listens Only)"
  }
  filter multiselect #fromQuestionFilter {
    optionsFrom: surveyDataset:TIME_OF_VISIT
    label: "Time of Visit (DN Listens Only)"
  }

  // filter reportingHierarchy #f_RestaurantHierarchy {
  //   reportingHierarchy: RestaurantHierarchy
  // }

  //AM filters

  filter multiselect #f_CaseStatus {
    optionsFrom: amTable:lk_3827
    label: "Case - Status"
  }
  filter multiselect #f_CaseCategories {
    optionsFrom: amTable:lk_3829
    label: "Case - Categories"
  }

  filter multiselect #f_CaseSeverity {
    optionsFrom: amTable:lk_3828
    label: "Case - Severity"
  }

  filter multiselect #f_CaseName {
    optionsFrom: amTable:CaseName
    label: "Case -  Trigger Names"
  }

//static filter is set but hidden
  filter singleselect #f_SurveyStatus {
    hide: false
    label: "Interview Status"

    option radio {
      label: "All Responses"
      value: _isnotnull(surveyDataset:status)
      //selected: true
    }

    option radio {
      label: "Completed interviews only"
      value: surveyDataset:status = "complete"

    }

    option radio {
      label: "Incomplete interviews only"
      value: surveyDataset:status = "incomplete"

    }
  } // end f_SurveyStatus
//this is to filter out test records. static filter is set but hidden
  filter singleselect #f_Production {
    hide: true
    label: "Production Interviews"
    option radio {
      label: "Production"
      value: _isnull(surveyDataset:test_resp) AND _isnull(surveyDataset.respondent:test_resp)
      selected: true
    }

    option radio {
      label: "Test"
      value: _isnotnull(surveyDataset.respondent:test_resp)

    }

  } // end f_Production
//static filter is set but hidden
  filter singleselect #f_HistoricalData {
    label: "Historical Data Filter"
    hide: true
    option radio {
      value: true
      label: "All Data"
      selected: true
    }
    option radio {
      value: _isnull(surveyDataset:hSMGData)
      label: "Current Data Only (no historical)"

    }
    option radio {
      value: _isnotnull(surveyDataset:hSMGData)
      label: "Historical Data Only"
    }


  } // end f_HistoricalData
  filter multiselect #f_Age {
    optionsFrom: surveyDataset:AGE
  }
  filter multiselect #f_Gender {
    optionsFrom: surveyDataset:GENDER
  }
  filter multiselect #f_Income {
    optionsFrom: surveyDataset:INCOME
  }

  filter multiselect #f_Region {
    optionsFrom: surveyDataset:RegionRecode
    label: "Region"
  }

} // end layoutArea toolbar
config pdfExport {
  pageSize: Letter
  pageOrientation: portrait, landscape
  pageScaling: fitToWidth
  exportMode: pdf
}

config report #reportConfig {
  logo: "/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/Logos/Delaware%20North%20site-logo.png"

  surveypid_kscvc: "p348419936952"
  surveypid_dnlistens: "p879777895877"
  surveypid_lodging: "p767600460264"
  surveypid_gaming: "p350899423091"
  surveypid_tours: "p195061967697"
  surveypid_lizard: "p895234707793"

  intvdate: surveyDataset:interview_start
  intvdate_ta: surveyDataset_TA:interview_start

  InvitedDate: .respondent:FirstEmailedDate
  CreatedDate: surveyDataset.respondent:CreatedDate

  //emailsSent: IN(.respondent:smtpStatus, "MessageSent", "Queued")
  emailsSent: count(.respondent:FirstEmailedDate) > 0

  //key metric fields
  nps_qid: surveyDataset:NPS
  osat_qid: surveyDataset:SAT
  value_qid: surveyDataset:Value

  //key metric fields
  nps_qid_ta: surveyDataset_TA:NPS
  osat_qid_ta: surveyDataset_TA:SAT
  value_qid_ta: surveyDataset_TA:Value

   //kpi targets 
  nps_target_score: 9

  //travel targets
  nps_travel_target: average(parseReal(SitesHierarchy:NPSTarget), SitesHierarchy:id = "DN_TRAVEL_HOSP")
  osat_travel_target: average(parseReal(SitesHierarchy:OSATTarget), SitesHierarchy:id = "DN_TRAVEL_HOSP")

  //lodging targets
  //nps_lodging_target: 46
  //osat_lodging_target: 53
  nps_lodging_target: average(parseReal(SitesHierarchy:NPSTarget), SitesHierarchy:id = "DN_PARKS")
  osat_lodging_target: average(parseReal(SitesHierarchy:OSATTarget), SitesHierarchy:id = "DN_PARKS")

  arrival_lodging_target: 61
  cleanliness_guestroom_lodging_target: 54
  cleanliness_bathroom_lodging_target: 54

  //gaming targets
  nps_gaming_target: average(parseReal(SitesHierarchy:NPSTarget), SitesHierarchy:id = "DN_GAMING")
  osat_gaming_target: average(parseReal(SitesHierarchy:OSATTarget), SitesHierarchy:id = "DN_GAMING")

  //KSCVC targets
  nps_kscvc_target: "TBD"
  //osat_kscvc_target: 70
  osat_kscvc_target: average(parseReal(SitesHierarchy:OSATTarget), SitesHierarchy:id = "1")

  //KSCVC targets
  nps_tours_target: "TBD"
  osat_tours_target: "TBD"

  restaurant_osat_target: 50

  nps_target: 61
  osat_target: 68
  ltc_target: 80
  promoters_target: 75
  problem_res_osat_target: 37

  sentiment_target_score: 2

  monthly_timeframe: "-12 month"

  suppressCriteriaMin: countif(surveyDataset:status = "complete") < 1
  KDAMinimumSampleSize: 10
  DNListensNonTravelLocations: "NFSP", "YGS", "BKT", "HHC", "JCW", "MRB", "TGB", "GGA", "SGB"
  DNListensParkLocations: "NFSP", "YGS"
  DNListensRestaurantLocations: "BKT", "HHC", "JCW", "MRB", "TGB", "GGA", "SGB"
  AustraliaLocations: "MBCR", "40765", "51906", "42458" //mindil, lizard, blacktown
  AustraliaPageLocations: "51906", "42458"  //lizard, blacktown
  ResponseRateNote: "NOTE: Response Rate = (# Respondents who answered NPS) / (# Invited)"

  HistoricalBenchmarksNote: "Threshhold for cell formatting = 4.00"
  PercentWithinCategoryNPS: "% within category: Promoters (9-10), Passives (7-8), Detractors (0-6)"
  PercentWithinCategory: "% within category: Top (4-5), Middle (3), Bottom (1-2)"

  aboveTargetLabel: "Above target"
  belowTargetLabel: "Below target"
  atTargetLabel: "At target"

  info_CardBackgroundColor: #F7F6D9
  selector_CardBackgroundColor: #F7F6D9

  nps_infoText: "The Net Promoter Score®, or NPS®, is a way of assessing the level of loyalty that a customer has toward an organization. We first ask a question about the customer's likelihood to recommend us:

ʺBased on your recent visit, on a scale from 0 to 10, how likely are you to recommend this location to a friend or family member? ʺ

Customers rating a 9 or 10 are called Promoters - these are the most favorable customers; on the other end of the spectrum, we have Detractors - those who rate from 0 to 6 on the scale. Customers rating 7 or 8 are put into a category called Passives.

To calculate the NPS®, we take the percentage of Promoters and subtract the percentage of Detractors. This means that NPS can fall on a scale between -100 (no Promoters) to 100 (all Promoters).

What should we do with this information? It can help with our efforts to act on customer insight - for example, Promoters are customers who are more likely to buy more (or different) products; they can also be great references. Detractors, on the other hand, often provide insight on areas of friction that we should consider Fixing."

  osat_infoText: "The overall satisfaction question assesses how happy the guest is with their entire experience with us. We also look at satisfaction on specific elements of their visit; these are reported separately. 

Satisfaction is measured on a five-point scale:

Very Dissatisfied
Somewhat Dissatisfied
Neither Dissatisfied Nor Satisfied
Somewhat Satisfied
Very Satisfied

Where a higher score is better.

We look at satisfaction based on the percentage of guests rating us as ʺVery Satisfiedʺ. We also report the average as well as the percentage who are dissatisfied (ʺSomewhat Dissatisfiedʺ or ʺVery Dissatisfiedʺ).

The satisfaction (OSAT) KPI gives us a sense for the holistic nature of their experience with their visit - this is the culmination of all the aspects of their interaction, which we drill into. OSAT gives us the ʺbig pictureʺ of the experience; to make it actionable, we need to break it down further (which our dashboards allow us to do easily)."

  value_infoText: "The overall value question assesses how guests evaluate the satisfaction of their experience relative to the amount of money spent. We often look at value on specific elements of their visit; these are reported separately. 

Value is measured on a five-point scale:

Poor Value
Marginal Value
Good Value
Very Good Value
Extremely Good Value

Where a higher score is better.

We look at value based on the percentage of guests rating us as an ʺExtremely Good Valueʺ or ʺVery Satisfied.ʺ 

The Value KPI gives us a sense for how guests view experience through an economic lens. Focusing on value instead of price alone is important, as guest will often accept higher prices when their satisfaction levels are at a commensurate level."



  kda_descriptionText: "This analysis looks for patterns in the data to identify how guest ratings on certain experiences influence their likelihood to recommend us to friends and family. This shows us where to target improvement initiatives at a strategic level."
  kda_quadrantColors_default: #ED1C24, #FFBD5B, #7A9A01, #00B2A9, #333333
  kda_quadrantColors: #ED1C24, #7A9A01, #FFBD5B, #00B2A9, #333333
  kda_quadrantTitles: "Fix First", "Leverage/Promote", "Consider Fixing", "Maintain/Monitor"
  kda_warningText: "* Item does not significantly add power to the analysis; please exercise caution when analyzing this variable."

  kda_infobox_label_correlation: "Key Driver Analysis (Correlation-Based)"
  kda_infobox_info_correlation: "**Correlation-Based Key Driver Analysis** is a statistical technique that shows the 1:1 relationship between individual aspects of the customer experience on a customer's overall satisfaction. This technique provides a framework for prioritizing action in a strategic manner. The analysis provides four outcomes:

1) ***Leverage/Promote*** - These are aspects that are important to customers that you perform well at; the strategy here is to maintain your current level of performance and promote these as differentiators.

2) ***Maintain/Monitor*** - These are things where you perform well, but are less important to customers at this time. These are areas that you should maintain at their current performance.

3) ***Fix First*** - These are areas that are important to customers, but your performance, relatively speaking, is weaker. These are the areas where improvements will generate the greatest lift from a customer sentiment perspective.

4) ***Consider Fixing*** - These are areas that, while your performance is weaker, are not areas of importance to customers. Focus on these areas after you have implemented improvements in the ***Fix First*** category.

Correlation-based analysis is not as robust as full regression-oriented analysis; however, it can be preferred when there is considerable skip patterns in data, as it allows for more cases to be included in the analysis than regression would.

It is important to note that Key Driver Analysis looks at the world as it is today - if something happens within your market (a disruptive product or service, or a new disruptive competitor, for example), then the underlying model that is being shown may change, and your drivers could change in terms of their impact."

  kda_infobox_label_regression: "Key Driver Analysis (Regression-Based)"
  kda_infobox_info_regression: "**Key Driver Analysis** is a statistical technique that shows the relationships among a series of aspects of the customer experience on a customer's overall satisfaction. This technique provides a framework for prioritizing action in a strategic manner. The analysis provides four outcomes:

1) ***Leverage/Promote*** - These are aspects that are important to customers that you perform well at; the strategy here is to maintain your current level of performance and promote these as differentiators.

2) ***Maintain/Monitor*** - These are things where you perform well, but are less important to customers at this time. These are areas that you should maintain at their current performance.

3) ***Fix First*** - These are areas that are important to customers, but your performance, relatively speaking, is weaker. These are the areas where improvements will generate the greatest lift from a customer sentiment perspective.

4) ***Consider Fixing*** - These are areas that, while your performance is weaker, are not areas of importance to customers. Focus on these areas after you have implemented improvements in the ***Fix First*** category.

It is important to note that Key Driver Analysis looks at the world as it is today - if something happens within your market (a disruptive product or service, or a new disruptive competitor, for example), then the underlying model that is being shown may change, and your drivers could change in terms of their impact."


//Palettes

  palette #multicolors1_palette {
    colors: #fa8072, #C7EA46, #104b6d, #7fffd4, #cec0b1, #737fc9, #C154C1, #cccccc, #F0E442, #155126,#7fffd4, #5310f0, #eac328, #82252a,#999999
    label: "Multi Colors 1 palette"
  }

  palette #multicolors2_palette {
    colors: #999999, #aee39a, #115e41, #4bc8e6, #40527a, #e9b4f5, #9d42b7, #78ee5a, #769d31, #21f0b6, #82252a, #fc7459, #6b4c33, #d18f60, #fd1e6e, #e9d737
    label: "Multi Colors 2 palette"
  }

  palette #redtogreen11ptscale {
    colors: #a50026, #d73027, #f46d43, #fdae61, #fee08b, #ffffbf, #d9ef8b, #a6d96a, #66bd63, #1a9850, #006837, #333333
  }


  palette #redtogreen5ptscale {
    colors: #d73027, #fdae61, #fee08b,  #a6d96a,  #1a9850,  #333333
  }

  palette #redtogreen3ptscale {
    colors: #d73027, #fdae61, #1a9850,  #333333
  }

  palette #redtogreen2ptscale {
    colors: #F3614D, #1a9850, #93949a
  }

  palette #greentored2ptscale {
    colors: #1a9850, #F3614D,  #333333
  }
  palette #copy_of_greentored2ptscale {
    colors: #1a9850, #93949a, #333333
    label: "2ptscale"
  }
  palette #copy_of_copy_of_greentored2ptscale {
    colors: #93949a, #1a9850, #333333
    label: "2ptscale reversed"
  }

  palette #kpi_palette {
    colors: #0096db, #58E2C0, #A75CD3, #000000
    label: "KPI colors palette"
  }


  palette #threecolor_palette {
   // colors: #98EE71,#FFBD5B,#F76473,#000000,#A6A6A6
    colors: #519B14, #FFBD5B, #FA5263, #000000

    label: "3 colors palette (reversed)"
  }

  palette #threecolor_palette_reversed {
    colors: #FA5263,#FFBD5B, #519B14, #000000
    label: "3 colors palette"
  }

  palette #nps_categories_palette {
    colors: #519B14, #FFBD5B, #FA5263, #000000
    label: "NPS Categories palette (reversed)"
  }

  palette #nps_palette_reversed {
    colors: #FA5263, #FFBD5B, #519B14, #000000
    label: "NPS Categories palette"
  }

  palette #nps_and_cats_palette {
    colors: #0096db, #FA5263,#FFBD5B, #519B14, #000000
    label: "NPS and Categories colors palette"
  }

  palette #survey_metrics_palette {
    colors: #0096db, #fdae61, #E85328, #000000
    label: "Survey Metrics palette"
  }



  palette #dot_palette {
    colors: #A4D65E
    label: "Dot palette"
  }
  palette #copy_of_dot_palette {
    colors: "#af5dd5"
    label: "Purple"
  }


//number formatters
  formatter number #oneDecimalFormatter {
    decimalSeparator: "."
    label: "oneDecimalFormatter"
    numberDecimals: 1
    integerSeparator: ","
    keepTrailingZeros: true
    shortForm: false
  }

  formatter number #noDecimalNumber {
    decimalSeparator: "."
    label: "noDecimalNumber"
    integerSeparator: ","
    numberDecimals: 0
  }

  formatter number #oneDecimalNumber {
    decimalSeparator: "."
    label: "oneDecimalNumber"
    integerSeparator: ","
    numberDecimals: 1
    keepTrailingZeros: true
  }

  formatter number #twoDecimalNumber {
    decimalSeparator: "."
    label: "twoDecimalNumber"
    integerSeparator: ","
    numberDecimals: 2
    keepTrailingZeros: true
  }

  formatter number #percentNumber {
    decimalSeparator: "."
    label: "percentNumber"
    postfix: "%"
    integerSeparator: ","
    numberDecimals: 0
    keepTrailingZeros: true
    shortForm: true
  }
  formatter number #noDecimalPercent {
    decimalSeparator: "."
    label: "noDecimalPercent"
    integerSeparator: ","
    postfix: "%"
    numberDecimals: 0
    //shortForm: true
  }

  formatter number #oneDecimalPercent {
    decimalSeparator: "."
    label: "oneDecimalPercent"
    integerSeparator: ","
    postfix: "%"
    keepTrailingZeros: false
    numberDecimals: 1
    //shortForm: true
  }

  formatter number #baseNumberFormatter {
    decimalSeparator: "."
    label: "noDecimalNumber"
    integerSeparator: ","
    numberDecimals: 0
    shortForm: false
    prefix: "(n = "
    postfix: ")"
  }

   //color formatters
  formatter color #neutral {
    thresholds: #848587 >= 0
    label: "neutral"
  }
  formatter color #positive {
    thresholds: #62B31C >= 0
    label: "positive"
  }
  formatter color #negative {
    thresholds: #D40001 >= 0
    label: "negative"
  }
  formatter color #colorFormatter {
    thresholds: #62B31C >= 9, #ff8e00 >= 7, #D40001 >= 0
    label: "backgroundColorFormatter2"
  }

  formatter color #dotColorFormatter {
    thresholds: #1D78BA >= 0
  }

  formatter color #percOfTotal {
    thresholds: #1D78BA >= 0%
    label: "percOfTotal"
  }

  formatter color #NPS_promoters {
    thresholds: #519B14 > 0
  }

  formatter color #NPS_passives {
    thresholds: #FFBD5B > 0
  }

  formatter color #NPS_detractors {
    thresholds: #FA5263 > 0
  }

  formatter color #openCasesColorFormatter_1 {
    label: "opencases"
    thresholds: #3DD864 >= 0
  }

  formatter color #closedCasesColorFormatter_1 {
    label: "closedcases"
    thresholds: #3b9cd8 >= 0
  }

  formatter color #inprogressCasesColorFormatter_1 {
    label: "inprogresscases"
    thresholds: #E7BC56 >= 0
  }

  formatter color #overdueCasesColorFormatter_1 {
    label: "overduecases"
    thresholds: #E96D25 >= 0
  }

  formatter color #TableBackgroundColorFormatter {
    label: "Red Amber Green Background (5 pt)"
    thresholds: #EEF7EA >= 5, #FFF5E7 >= 3, #FFECEE < 3
  }
  formatter color #copy_of_TableBackgroundColorFormatter {
    label: "Red Amber Green Background (NPS)"
    thresholds: #EEF7EA >= 50, #FFF5E7 >= 0, #FFECEE < 0
  }

  formatter color #background_diff_goal {
    thresholds: #A52B31 <= -20, #DA6F74 <= -10, #72BF44 >= 20, #AAD98F >= 10
    label: "background_diff_goal"
  }
  formatter color #text_diff_goal {
    thresholds: #ffffff <= -20, #000000 <= -10, #000000 >= 20, #000000 >= 10
    label: "text_diff_goal"
  }

  formatter color #background_diff_previous {
    thresholds: #A52B31 <= -20, #DA6F74 <= -10, #72BF44 >= 20, #AAD98F >= 10
    label: "background_diff_previous"
  }
  formatter color #text_diff_previous {
    thresholds: #ffffff <= -20, #000000 <= -10, #000000 >= 20, #000000 >= 10
    label: "text_diff_previous"
  }

  formatter color #background_zeros_formatter {
    thresholds: #DA6F74 < 1
    label: "background_zeros_formatter"
  }
  formatter color #text_zeros_formatter {
    thresholds: #000000 >= 0
    label: "text_zeros_formatter"
  }

//date formatters
  formatter date #monthShort {
    inputFormat: YYYYMM
    formatString: "MMM YYYY"
  }

  formatter date #month {
    inputFormat: YYYYMM
    formatString: "MMMM YYYY"
  }
  formatter date #quarter {
    inputFormat: YYYYQQ
    //formatString: "\Q\t\r Q YYYY"
    formatString: "YYYY \Q\t\r Q"
  }

  formatter date #week {
    inputFormat: YYYYWW
    formatString: "\W\e\e\k W YYYY"
  }

  formatter date #dateFormatDay {
    inputFormat: "YYYYMMDD"      //put the current format of how the date comes out on the chart here
    formatString: "MM-DD-YYYY"  //use a slash to include text within the date format
  }


//TA formatters
  formatter color #sentimentindicator {
    thresholds: #98EE71  >=1, #fee090 >-1, rgba(244, 88, 88, 0.867) <= -1
    defaultValue: transparent
  }
  formatter color #sentimentindicatortext {
    thresholds: #333333 >=1, #333333 >-1, #FFFFFF <=-1
    defaultValue: transparent
  }
  formatter color #copy_of_sentimentindicatortext {
    thresholds: #333333 >= 50, #333333 >= 0, #333333 < 0
    defaultValue: transparent
    label: "Text (NPS)"
  }
  formatter color #sentimentindicator2a {
    thresholds: transparent >= 0
  }

  formatter color #sentimentindicator2text {
    thresholds: #508F19  >= 3, #848587 >=2, #D40001 >=1
  }
  formatter color #sentimentindicatortextValue2 {
    thresholds: Positive >= 3, Neutral >= 2, Negative >=1, None<0
    label: "Sentiment Indicator Text"
  }

  formatter color #sentimentindicatortext2 {
    thresholds: #333333 >= 3, #333333 >= 2, #FFFFFF >=1
    //thresholds: #333333 >= 0.25, #333333 >= -0.25, #FFFFFF >= -5
  }

  formatter color #sentimentindicator2 {
    thresholds: #98EE71 >= 3, #fee090 >=2, #F45858 >=1
    //#e8f8e0 comments lighter green
    //thresholds: #8BCB24 >= 0.25, #fee090 >= -0.25, #F45858 >= -5
  }



  formatter color #sentimentindicator1 {
    thresholds: #6DC548 >= 9, #FFC832 >= 7, #F3614D >= 0, #F9F9F9 < 0
    defaultValue: transparent
  }
  formatter color #sentimentindicator1text {
    thresholds: #000000 >= 9, #000000 >= 7, #000000 >= 0, #F9F9F9 < 0
    defaultValue: transparent
  }

  formatter color #sentimentindicator_bg_5pt {
    thresholds: #6DC548 >= 4, #FFC832 >= 3, #F3614D >= 0, #F9F9F9 < 0
    defaultValue: transparent
  }
  formatter color #sentimentindicator_text_5pt {
    thresholds: #000000 >= 4, #000000 >= 3, #000000 >= 0, #F9F9F9 < 0
    defaultValue: transparent
  }

  formatter color #npssegmentindicator2 {
    thresholds: #8BCB24 >= 3, #fee090 >=2, #F45858 >=1
  }
  formatter color #npssegmentindicatortext2 {
    thresholds: #FFFFFF >= 3, #333333 >= 2, #FFFFFF >=1
  }
  formatter color #npssegmentindicatortextValue2 {
    thresholds: Promoter >= 3, Passive >= 2, Detractor >=1,None<0
  }

  palette answerList #paletteNegNeuPos {
    item {
      code: "Negative"
      color: #F76473
    }
    item {
      code: "Neutral"
      color: #FFBD5B
    }
    item {
      code: "Positive"
      color: #98EE71
    }
  }

  palette #palettePosNegNueReverse {
    colors: #98EE71,#FFBD5B,#F76473,#000000,#A6A6A6
    label: "palette Pos Neg Nue Reverse"
  }

  //TA COLOR FORMATTERS
  formatter color #colorPositive {
    label: "Positive"
    thresholds: #519B14 >= 0
  }
  formatter color #colorNeutral {
    label: "Neutral"
    thresholds: #FFBD5B >= 0
  }
  formatter color #colorNegative {
    label: "Negative"
    thresholds: #FA5263 >= 0
  }
  formatter color #sentimentIndicatorWording {
    label: "Sentiment Indicator Wording"
    //thresholds: Positive > 0, Neutral = 0, Negative < 0
    thresholds: Positive >= 3, Neutral >= 2, Negative >=1,None<0
  }

  formatter color #dropOffDefaultFormatter {
    label: "One Color"
    thresholds: #004d63 >= 0, #004d63 < 0
    // This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter color #taSentimentColorDefaultFormatter {
    label: "TA Sentiment Numeric Background"
    thresholds: #98EE71 > 0.25, #fee090 >= -0.25, #F56E6E >= -5
    // This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter color #copy_of_taSentimentColorDefaultFormatter {
    label: "Copy of TA Sentiment Numeric Background"
    thresholds: #EEF7EA > 0.25, #FFF5E7 >= -0.25, #FFECEE >= -5
    // This default formatter was added to CDL when it was overridden in the widget library
  }

  formatter color #scoreNPS_green {
    thresholds: #98EE71 > 0
  }

  formatter color #scoreNPS_orange {
    thresholds: #FFBD5B > 0
  }

  formatter color #scoreNPS_red {
    thresholds: #F76473 > 0
  }

  formatter color #scoreNPS_grey {
    thresholds: #bdbcbc > 0
  }

  formatter color #scoreNPS_blue {
    thresholds: #7dbce3 > 0
  }

//target formatters for infographics
  formatter color #OverallOSATFormatter {
    thresholds: #62B31C >= 61, #E85328 < 61
  }

  formatter color #PromotersFormatter {
    thresholds: #62B31C >=67, #E85328 < 67
  }


  formatter color #gridDefaultBackgroundColorFormatter {
    label: "Red Amber Green Background"
    thresholds: #EEF7EA >= 95%, #FFF5E7 >= 90%, #FFECEE < 90%
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter color #gridDefaultValueColorFormatter {
    label: "Red Amber Green Percent (Grid)"
    thresholds: #388E3C >= 95%, #FF8E00 >= 90%, #D40000 < 90%
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter color #kpiColorDefaultFormatter {
    label: "Red Amber Green Percent (KPI)"
    thresholds: #62B31C >= 100%, #FF8E00 >= 80%, #D40001 < 80%
    defaultValue: "#007DB8"
// This default formatter was added to CDL when it was overridden in the widget library
  }
} // config reportConfig
page #page_MainOverview {
  label: "Executive Overview"
  access rules {
    rule claim {
      name: "UserSegment"
      //value: "All", "Travel"
      value: "Test"
    }
  }
  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }


  widget headline #headlineWidget_7 {
    label: "Delaware North Customer Listening Dashboard"

    size: large

    tile markdown #markdownTile_2 {
      value: "# Executive  Overview 
### This dashboard provides an overview of guests’ feedback about their experiences with our organization across Parks, Gaming, and THS. 
Data is collected through our Voice of Guest surveys, which are either deployed post visit or displayed through a QR code onsite. 

 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key Drivers that impact guest experience
- Trends
- A view of each property’s performance against their KPI goal
- Verbatims comments from guests
 
You can click on the filter icon in the upper left hand corner of the report to refine who is included in the report, including narrowing your focus to a single survey type. 
When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing).***
"

    }
    // tile button #buttonTile {
    //   value: "Go To Action Management"
    //   navigateTo: "page_CasesOverview"
    //   navigateOptions: "same_tab"
    //   //navigateFilter: surveyDataset:filterMeasure_DNListensTravelOnly()
    // }

  }
  widget kpi #kpiWidget_4 {
    label: "Parks Lodging OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    filter expression {
      value: surveyDataset:filterMeasure_LodgingSurvey()
      label: "Lodging Only"
    }


    // filter expression  {
    //   value: surveyDataset:filterMeasure_ExcludeAustraliaLocations()
    //   label: "Exclude Australia locations"
    // }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_lodging_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all lodging locations with Parks & Resorts.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_5 {
    label: "KSCVC OSAT"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    filter expression {
      value: surveyDataset:filterMeasure_KSCVCSurvey()
      label: "KSCVC Only"
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_kscvc_target
//target: average(parseReal(SitesHierarchySimplified:OSATTarget), SitesHierarchySimplified:id="1")
    }


    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **Kennedy Space Center Visitors Complex.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  } // end widget
  widget kpi #kpiWidget_6 {
    label: "Tours OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    filter expression {
      value: surveyDataset:filterMeasure_ToursSurvey()
      label: "Tours Only"
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_tours_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Tours.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_7 {
    label: "Gaming NPS®"
    size: small
    ignoreFilters: f_Location

    filter expression {
      value: surveyDataset:filterMeasure_GamingSurvey()
      label: "Gaming Only"
    }

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_ExcludeAustraliaLocations()
      label: "Exclude Australia locations"
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_gaming_target
    }
    infobox #infobox {
      label: "NPS®"
      info: "The Net Promoter Score®, or NPS®, is a way of assessing the level of loyalty that a customer has toward an organization. We first ask a question about the customer's likelihood to recommend us:

ʺBased on your recent visit, on a scale from 0 to 10, how likely are you to recommend this location to a friend or family member? ʺ

Customers rating a 9 or 10 are called Promoters - these are the most favorable customers; on the other end of the spectrum, we have Detractors - those who rate from 0 to 6 on the scale. Customers rating 7 or 8 are put into a category called Passives.

To calculate the NPS®, we take the percentage of Promoters and subtract the percentage of Detractors. This means that NPS can fall on a scale between -100 (no Promoters) to 100 (all Promoters).

What should we do with this information? It can help with our efforts to act on customer insight - for example, Promoters are customers who are more likely to buy more (or different) products; they can also be great references. Detractors, on the other hand, often provide insight on areas of friction that we should consider Fixing."
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all Gaming locations.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above.

Note: Australia locations have been excluded on this widget."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }

  }
  widget kpi #kpiWidget_8 {
    label: "Travel Hospitality NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    filter expression {
      value: surveyDataset:filterMeasure_DNListensTravelOnly()
      label: "DN Listens-Travel locations only"
    }

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all Travel Hospitality locations.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_9 {
    label: "Patina OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    filter expression {
      value: surveyDataset:filterMeasure_DNListensRestaurants()
      label: "DN Listens-Restaurant locations"
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.osat_travel_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Patina locations.**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_10 {
    label: "Australia Lodging NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_AustraliaLocations()
      label: "Australia Locations"
    }

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
     // target: @reportConfig.nps_lodging_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **All Australia lodging locations within Parks & Resorts.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget headline #headlineWidget_8 {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Exec_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget dataGrid #dataGridWidget_2 {
    label: "Parks - Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "This view displays a breakdown of the performance of all locations on our key performance indicators. This provides insight on how locations perform in a relative context.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_lodging), SitesHierarchySimplified:^hierarchy) > 0 OR count(:, selected(:survey_pid, @reportConfig.surveypid_kscvc), SitesHierarchySimplified:^hierarchy) > 0 OR count(:, selected(:survey_pid, @reportConfig.surveypid_tours), SitesHierarchySimplified:^hierarchy) > 0

    }

    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_current_counts {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        navigateTo: page_LodgingResponses

      }

    }

    column #column_current_NPS {

      label: "NPS®"

      // scope reportingPeriod {
      //   period: Current
      // }
      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        navigateTo: page_LodgingResponses
       // view: comparativeStatisticView
      }
    }

    column cut #column_Promoters {
      //value: recode(@reportConfig.nps_qid, @NPScats)
      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_LodgingResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    // column #NPSPosNegNeutral {
    //   label: " % within NPS® category "

    //   cell microchart {
    //     value: count(surveyDataset:)
    //     format: noDecimalNumber
    //           //extraValue: count(@reportConfig.nps_qid)
    //     breakdownBy cut {
    //       value: surveyDataset:NPSVal

    //      // value: LoyaltyGrid:value
    //     }
    //     microchart stacked100PercentBar {
    //       valuePosition: none
    //       palette: nps_palette_reversed
    //       notAnswered: false
    //       showTooltip: true
    //       percentFormat: oneDecimalPercent

    //     }
    //   }
    // }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Exec_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Lodging_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Exec_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_current_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_LodgingResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }

    column #column_OSATGoal {

      label: "OSAT Goal"

      format: noDecimalNumber

      cell {

        value: parseReal(SitesHierarchySimplified:OSATTarget)
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_OSAT_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_OSAT
        other: column_OSATGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Exec_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Lodging_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Exec_Timeframe_Selector.selected.selectBreakdownBy
        }

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget dataGrid #dataGridWidget_3 {
    label: "Gaming - Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "### This view displays a breakdown of the performance of all locations on our key performance indicators. This provides insight on how locations perform in a relative context.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }


    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_gaming), SitesHierarchySimplified:^hierarchy) > 0

    }

    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_current_counts {
      label: "n"
      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }

    }

    column #column_current_NPS {

      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        navigateTo: page_GamingResponses
       // view: comparativeStatisticView
      }
    }

    column #column_NPSGoal {

      label: "NPS® Goal"

      format: noDecimalNumber
      // scope reportingPeriod {
      //   period: Current
      // }
      cell {
        //for any locaitons without a target, set target to "TBD" in the table
        value: parseReal(SitesHierarchySimplified:NPSTarget)

        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_NPS_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_NPS
        other: column_NPSGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column cut #column_Promoters {
      //value: recode(@reportConfig.nps_qid, @NPScats)
      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_GamingResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }


    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column {
      label: "NPS® Trends" + " - " + @Exec_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Locations_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Exec_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_current_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_GamingResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }

    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Exec_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Locations_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Exec_Timeframe_Selector.selected.selectBreakdownBy
        }

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget dataGrid #dataGridWidget_6 {
    label: "Travel Hospitality - Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }
    // filter expression {
    //   value: depth(SitesHierarchySimplified:^hierarchy) >= 1
    // }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_dnlistens), SitesHierarchySimplified:^hierarchy) > 0

    }
    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row selectedFlat #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      labelStyle: nodeOnly
    //showTotal: true
    }

    column #column_current_counts {
      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
      }

    }

    column #column_current_NPS {
      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
       // target: parseReal(SitesHierarchy:NPSTarget)
        navigateTo: page_DNListensResponses
       //view: comparativeStatisticView
      }
    }

    column #column_NPSGoal {

      label: "NPS® Goal"

      format: noDecimalNumber

      cell {
        value: parseReal(SitesHierarchySimplified:NPSTarget)
        //value: average(numeric(Goals_CustomTable:nps_target))
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_NPS_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_NPS
        other: column_NPSGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column cut #column_Promoters {

      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_DNListensResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Exec_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Exec_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_DNListensResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }
    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Exec_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Exec_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

      }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget table #tableWidget {
    label: "Visitor Comments"
    size: "large"
    table: surveyDataset:

    showHeader: true
    sortOrder: descending
    sortColumn: comments

    headerNumberOfLines: 3
    stretchColumns: true

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000


    navigateTo: page_Indiv_Survey_Response
    description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response."


    select #OpenEnd_selector {
      label: "Select Question"
      options: item {
        label: "Visit Comments"
        value:  {
          selectQuestion: surveyDataset:VISIT_COMMENTS
          selectFilter: surveyDataset:VISIT_COMMENTS != ""
        }

      },
	    item {
        label: "Lodging Comments"
        value:  {
          selectQuestion: surveyDataset:LODGING_COMMENTS
          selectFilter: surveyDataset:LODGING_COMMENTS != ""
        }

      },
	    item {
        label: "Restaurant/Buffet Comments"
        value:  {
          selectQuestion: surveyDataset:RESTAURANT_COMMENTS
          selectFilter: surveyDataset:RESTAURANT_COMMENTS != ""
        }

      },
      item {
        label: "Problem Details"
        value:  {
          selectQuestion: surveyDataset:PROBLEM_DETAIL
          selectFilter: surveyDataset:PROBLEM_DETAIL != ""
        }

      },
      item {
        label: "Team Recognition"
        value:  {
          selectQuestion: surveyDataset:RECOG_DETAIL
          selectFilter: surveyDataset:RECOG_DETAIL != ""
        }

      }    

    } // end OpenEnd_selector
    filter expression {
      value: @OpenEnd_selector.selected.selectFilter
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }


    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }


    column response #comments {
      //sortBy: comment
      header: "Location: " + surveyDataset:LocationName
      footer: @reportConfig.intvdate
     // width: 300px
      enableColumnFilter: true
      comment: @OpenEnd_selector.selected.selectQuestion

    }


    // column value #SurveyName {
    //   label: "Survey"
    //   value: surveyDataset:survey_name
    //   enableColumnFilter: true
    //   align: center
    //   width: 150px

    // }


    column value #SurveyName {
      label: "Survey Name"
      value: surveyDataset:survey_name
      //value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 100px
    }

    column value #LocationName {
      label: "Location"
      value: demote(SitesHierarchy:language_text, surveyDataset:)
      //value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 200px
    }

    // column value #LoyaltyTier {
    //   label: "Loyalty Tier"
    //   value: surveyDataset:rank_description
    //   //value: surveyDataset:LocationName
    //   enableColumnFilter: true
    //   //value: surveyDataset:SitesHierarchy
    //   width: 100px
    // }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Rec"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    column metric #copy_of_metricColumn {
      label: "OSAT"
      value: score(@reportConfig.osat_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

  } // end widget
  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
} // end page
page #page_TravelOverview {
  label: "Travel Hospitality"

  access rules {
    rule claim {
      name: "UserSegment"
      value: "All", "Travel"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }

  filter expression {
    value: surveyDataset:filterMeasure_DNListensTravelOnly()
    label: "DN Listens-Travel locations only"
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  widget headline #headlineWidget_4 {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Travel Hospitality - Airports 
### This dashboard compiles survey data collected within airports through QR code surveys. This survey was previously referred to as the DN Listens survey. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatims comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a single airport. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }


    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_DNListensTravelOnly()
    }


    label: "Voice of Guest Dashboard"
  }


  widget kpi #kpiWidget_Overall_NPS {
    label: "Overall Subsidiary NPS®"
    size: small
    ignoreFilters: f_Location
    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all Travel Hospitality locations.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Overall Subsidiary OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.osat_travel_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Travel Hospitality locations.**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Travel Hospitality location(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Travel Hospitality location(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  }
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: oneDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: primary
      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
    }
  }
  widget headline #headlineWidget_totalOpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small

    //     tile text #textTile0 {
    //   value: "" + @currentUser.Node
    //   fontSize: 20
    // }

    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_Recognize {
    label: "Recognize a Team Member?"
    hide: true

    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"


    category cut #cutCategory {
      value: :PROBLEM

    }
    palette: redtogreen2ptscale
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  }
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Travel_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Travel_Timeframe_Selector.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Travel_Timeframe_Selector.selected.selectFilter
    // }


    // select #OSAT_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_7 {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
#### **Goals shown are current year 2024 goals; please keep this in mind if you change the reporting period.**
[Click here to open the pdf 'THS Annual NPS Goals Review'](/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/goals/DelawareNorth_THS_Annual_Goals.pdf)
"


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }
    // filter expression {
    //   value: depth(SitesHierarchySimplified:^hierarchy) >= 1
    // }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_dnlistens), SitesHierarchySimplified:^hierarchy) > 0

    }
    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row selectedFlat #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      labelStyle: nodeOnly
    //showTotal: true
    }

    column #column_current_counts {
      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
      }

    }

    column #column_current_NPS {
      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
       // target: parseReal(SitesHierarchy:NPSTarget)
        navigateTo: page_DNListensResponses
       //view: comparativeStatisticView
      }
    }

    column #column_NPSGoal {

      label: "NPS® Goal"

      format: noDecimalNumber

      cell {
        value: parseReal(SitesHierarchySimplified:NPSTarget)
        //value: average(numeric(Goals_CustomTable:nps_target))
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_NPS_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_NPS
        other: column_NPSGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column cut #column_Promoters {

      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_DNListensResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_DNListensResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }
    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

      }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. 
[THS Annual NPS Goals Review](/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/goals/DelawareNorth_THS_Annual_Goals.pdf)"
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

    fixedHeader: true
  } // end widget
  widget keyDrivers #keyDriversWidget_OSAT_Travel {
    label: "What Drives Guest Satisfaction?"
    algorithm: regression
    dependentVariable: @reportConfig.osat_qid
    independentVariables: surveyDataset:SAT_DRIVERS.quality, surveyDataset:SAT_DRIVERS.value, surveyDataset:SAT_DRIVERS.variety, surveyDataset:SAT_DRIVERS.speed, surveyDataset:SAT_DRIVERS.staff
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    quadrantColors: @reportConfig.kda_quadrantColors
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression
    }
    description: "This analysis looks for patterns in the data to determine how guest ratings on certain experiences influence their overall satisfaction with their visit. This shows us where to target improvement initiatives."
    importanceLimit: 0.2
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_OSAT_Travel
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments with Text Analytics**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  }
  widget comments #commentsWidget_Dining {
    label: "Comments with Text Analytics sentiment and categories"
    size: large
    table: textAnalyticsDataset_Dining.overallScore:
    sortOrder: descending
    sortColumn: responseColumn

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000
    navigateTo: page_Indiv_Survey_Response_TA

    infobox #infobox {
      label: "Information"
      info: "This widget shows all verbatim comments, and the comment's overall sentiment or other contextual variables related to the comment. 
- Overall sentiment is measured for all the text in a comment field rather than parts of it.
- Overall sentiment ranges from -5 to 5. 0 is neutral or mixed. 
- Tags under each comment represent the topic categories associated with this comment. Tags are color-coded red for negative, yellow for neutral/mixed and green for positive. 
- Columns are filterable.
- Clicking anywhere on a comment will bring you to the Response-level results."
    }


    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: large
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: large
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
    }

    group question #questionGroup {
      label: "All Comments"
      comment: textAnalyticsDataset_Dining.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Dining.overallScore:text != ""
      }
    }
    column response #responseColumn {
      sortBy: footer
      //header: "Claim #" + surveyDataset:ClaimNbr
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta

      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "Comment Field"
      value: textAnalyticsDataset_Dining.overallScore:variable
      enableColumnFilter: true
      width: 150px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #StoreName {
      label: "Store / Restaurant"
      value: surveyDataset_TA:STORE_INFO
      enableColumnFilter: true
      //value: surveyDataset_TA:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Dining:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Dining:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 125px
    }

    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    column metric #metricColumn_NPS {
      label: "NPS"
      value: score(@reportConfig.nps_qid_ta)
      enableColumnFilter: true
      //filterable: true
      width: 125px
      align: center
      view: colorcoding
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_OSAT {
      label: "SAT"
      value: score(@reportConfig.osat_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }


    description: "**Note: To filter on Overall Sentiment, enter 3 for Positive, 2 for Neutral, 1 for Negative**
    **Note: To filter on NPS Segment, enter 3 for Promoters, 2 for Passives, 1 for Detractors**"


  } // end widget
  widget chart #TopTopics_chartWidget {

  //  label: @TANumTopics_Selector.selectedLabel + " " + @TACategoryLevels_Selector.selectedLabel + " by Volume"
    label: "Top 10 Text Analytics Topics by Volume"

    size: large
    animation: false
    gridLines: false
    legend: bottomCenter
    layout: "horizontal"
    palette: palettePosNegNueReverse

    hide: false

    filter expression {
      //value: depth(textAnalyticsDataset_Dining.model:^parent) = @TACategoryLevels_Selector.selected
      value: depth(textAnalyticsDataset_Dining.model:^parent) = 1
    }

    series #volume1 {
      label: "Mentions"
      value: textAnalyticsDataset_Dining:categoryCountTASet1()
      format: noDecimalNumber
      //navigateFilter: some(textAnalyticsDataset_Dining.categoryScore:, true, textAnalyticsDataset_Dining.categoryScore:)
      //navigateTo: dd_CategoryResultsByThemeComments
      navigateTo: dd_SentimentComments_Dining

      breakdownBy cut {
        value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      }
      percent: false
      chart bar {
        mode: stacked
        maxBarSize: 65
      }
    }
    category selectedFlat {
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
     // takeTop: @TANumTopics_Selector.selected
      takeTop: 10
      sortBy: "volume1"
      sortOrder: descending
    }


    axis secondary {
      label: "Category Sentiment"
      hide: true
    }

    axis category #categoryAxis {

      textSize: 150
      orientation: "-45"
    }
    axis primary {
      format: noDecimalNumber
    }
    navigateTo: "page_Parks_Overview"
  } // end widget
  // widget headline #headlineWidget_8 {
  //   label: "Text Analytics Sentiment Trends"
  //   size: large
  //   cardBackground: @reportConfig.selector_CardBackgroundColor


  //   select #TA_Timeframe_Selector_Dining {
  //     label: "Select a Timeframe"
  //     options: @valueSet_date_ranges.items

  //   } // end selector
  //   tile markdown #markdownTile {
  //     value: "### The section displays sentiment trends."
  //   }

  // } // end widget
  widget chart #SentimentTrends_chartWidget {
    label: "Text Analytics Sentiment Components Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    size: large
    animation: true
    gridLines: horizontal
    legend: bottomCenter
    removeEmptyCategories: true
    //navigateTo: dd_SentimentComments
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Timeframe_SelectorTA1.selected.selectFilter
    // }

    infobox #infobox {
      label: "Information"
      info: "This widget shows the % distribution of overall sentiment over time. Time period break (first drop-down menu) and sentiment group base (second drop-down menu) may be selected. The distribution of the sentiment group is based on either respondents or comments for (All, positive, neutral/mixed, or negative). 
- Overall sentiment is measured for all the text in a comment field rather than parts of it. 
- Hover over the dots for more info.
- Clicking on a bar or dot will take you to the category results for that time period."
    }

    series #series_primary {
      chart bar {
        mode: "stacked100Percent"
        dataLabel: percentThenValue
        barSize: 75
        maxBarSize: 75
      }
      value: textAnalyticsDataset_Dining:overallResponseBaseTASet1()
      label: "% distribution of respondents by sentiment group"
      format: noDecimalNumber
     // format: @metric_selector.selected.cellFormat
      palette: paletteNegNeuPos
      navigateTo: dd_SentimentComments_Dining

      breakdownBy cut #cutBreakdownby {
        value: textAnalyticsDataset_Dining:responseSentimentGroup()
      }
    }

    series #series_secondary {
      value: textAnalyticsDataset_Dining:overallAverageTASet1()
      format: oneDecimalNumber
      label: "Average Sentiment"
      isSecondary: true
      chart line {
        lineWidth: 3
        dotSize: 7
        dotColorFormat: taSentimentColorDefaultFormatter
        connectNulls: true
        showDotValue: true
      }
      palette: palettePosNegNueReverse
    }


    category date #cutByDate {
      value: @reportConfig.intvdate_ta
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

    }

    chartMargin {
      top: 20
    }
    axis primary {
      label: "%"
      format: percentNoDecimal
      minValue: 0
      maxValue: 100
    }
    axis category {
      orientation: -45
      textSize: 75
    }
    axis secondary #secondaryAxis {
      label: "Sentiment (-5 to 5)"
      minValue: -5
      maxValue: 5
      format: noDecimalNumber
    }
    base {
      value: textAnalyticsDataset_Dining:overallResponseBaseTASet1()
      format: baseNumberFormatter
    }
    removeEmptySeries: true
  } // end widget
  widget headline #CatsAndSentiment_headlineWidget {
    label: "Text Analytics Categories & Sentiment Analysis"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #HierView_Selector {
      label: "Select a View"
      options: @valueSet_hierarchy_views.items

    } // end selector
    tile markdown #markdownTile {
      value: "###"
    }

  } // end widget
  widget dataGrid #CatsAndSentiment_HierView {
    label: "Text Analytics Categories & Sentiment - Hierarchical View"
    size: "large"

    hide: @HierView_Selector.selected != 1

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedHierarchy #comparisonRow {
      sortBy: "/percentTotalComments"
      sortOrder: descending
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:percentageOfCommentsTASet1()
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Dining:categoryCountTASet1()
        format: noDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

        }
        format: oneDecimalNumber

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Dining:categoryCount()
        extraValue: textAnalyticsDataset_Dining:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
  widget dataGrid #CatsAndSentiment_FlatView {
    label: "Text Analytics Categories & Sentiment - Flat view"
    size: "large"
    //navigateTo: dd_CategoryResultsByThemeComments

    hide: @HierView_Selector.selected != 2

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector


    row selectedFlat #comparisonRow {
      sortOrder: descending
      sortBy: "/percentTotalComments"
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:percentageOfCommentsTASet1()
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Dining:categoryCountTASet1()
        format: noDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Microcharts_Timeframe_Selector.selected.selectFilter
      // }
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()

        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

        }
        format: oneDecimalNumber

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Dining:categoryCount()
        extraValue: textAnalyticsDataset_Dining:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }

    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }
  } // end widget
  widget table #tableWidget_Comments_Hist {
    label: "Historical Comments (SMG)"
    size: "large"
    table: surveyDataset:

    showHeader: true
    sortOrder: descending
    sortColumn: comments

    headerNumberOfLines: 3
    stretchColumns: true

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response
    description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response.

Note: ʺReason for Recommendationʺ was added in the survey starting February 6, 2023. ʺTell us about your Experienceʺ was asked prior to that and continued until Apr 27, 2023."

    select #histOpenEnd_selector {
      label: "Select Question"
      options: item {
        label: "Reason for Recommendation"
        value:  {
          selectQuestion: surveyDataset:SMG_RecmdComments
          selectFilter: surveyDataset:SMG_RecmdComments != ""
        }

      },
	    item {
        label: "Tell us about your Experience"
        value:  {
          selectQuestion: surveyDataset:SMG_ExpComments
          selectFilter: surveyDataset:SMG_ExpComments != ""
        }

      }
    } // end histOpenEnd_selector
    filter expression {
      value: @histOpenEnd_selector.selected.selectFilter
    }
    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }


    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }


    column response #comments {
      //sortBy: comment
      header: "Location: " + surveyDataset:LocationName
      footer: @reportConfig.intvdate
     // width: 300px
      enableColumnFilter: true
      comment: @histOpenEnd_selector.selected.selectQuestion

    }

    column value #LocationName {
      label: "Location"
      value: demote(SitesHierarchy:language_text, surveyDataset:)
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #StoreName {
      label: "Store / Restaurant"
      value: surveyDataset:STORE_INFO
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Recm'd"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    // column metric #copy_of_metricColumn {
    //   label: "OSAT"
    //   value: score(@reportConfig.osat_qid)
    //   enableColumnFilter: true
    //   width: 100px
    //   align: center
    //   view: colorcoding_5pt

    // }

  } // end widget
  widget markdown #markdownWidget_PerformanceTrends {
    markdown: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    size: large
  }
  widget dataGrid #dataGridWidget_SatDrivers {
    label: "Satisfaction Drivers"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_DRIVERS$field
      total: none

    }
    column #column_current_counts {
      value: count(:SAT_DRIVERS$value)
      label: "Number of Responses"
      cell {
        value: count(:SAT_DRIVERS$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

    description: "Note: Variety and Value measures included in survey starting April 27, 2023.  Quality, Speed of Service, and Friendliness of Staff were included in the survey starting February 6, 2023.

Note: 'N/A' responses have been filtered out of the results below."
  } //end widget
  widget dataGrid #dataGridWidget_Sat_TimeOfDay {
    label: "Satisfaction By Time of Day"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    // sort rows {
    //   sortBy: "/Satisfaction"
    //   sortOrder: descending
    // }

    row cut {
      value: surveyDataset:TIME_OF_VISIT
      total: none

    }
    column #column_current_counts {
      value: count(surveyDataset:TIME_OF_VISIT)
      label: "Number of Responses"
      cell {
        value: count(surveyDataset:TIME_OF_VISIT)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }


    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023"
  } //end widget
  widget chart #dataGridWidget_Sat_TimeOfVisit {
    label: "Satisfaction By Time of Visit" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: multicolors1_palette
   // ignoreFilters: reportingPeriodFilter

    // select #TimeofDay_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 75
      right: 25
    }

    series #series {
      chart line {
        showDotValue: false

      }

      value: top1percent(@reportConfig.osat_qid)
      format: oneDecimalPercent

      isSecondary: false
      breakdownBy cut {
        value: surveyDataset:TIME_OF_VISIT

      }
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }


    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "% Very Satisfied"
      minValue: 50
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }


    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
  } // end widget
} // end page
page #page_RestaurantsOverview {
  label: "Restaurants"

  access rules {
    rule claim {
      name: "UserSegment"
      //value: "All", "Travel"
      value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }

  filter expression {
    value: surveyDataset:filterMeasure_DNListensRestaurants()
    label: "DN Listens-Restaurant locations"
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  widget headline #headlineWidget_4 {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Restaurants: Patina & Sportservice
### This dashboard compiles survey data collected within Patina and Sportservice Restaurants, collected through QR code surveys. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Trends
- Verbatims comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a single airport. 
When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }


    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_DNListensNonTravel()
    }


    label: "Voice of Guest Dashboard"
  }


  widget kpi #kpiWidget_Overall_NPS {
    label: "Restaurant NPS®"
    size: small
    ignoreFilters: f_Location
    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all Restaurant locations.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Restaurant OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.osat_travel_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Restaurant locations.**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Restaurant location(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Restaurant location(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  }
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: oneDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: primary
      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
    }
  }
  widget headline #headlineWidget_totalOpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small

    //     tile text #textTile0 {
    //   value: "" + @currentUser.Node
    //   fontSize: 20
    // }

    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_Recognize {
    label: "Recognize a Team Member?"
    hide: true

    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"


    category cut #cutCategory {
      value: :PROBLEM

    }
    palette: redtogreen2ptscale
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  }
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Travel_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Travel_Timeframe_Selector.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Travel_Timeframe_Selector.selected.selectFilter
    // }


    // select #OSAT_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }
    // filter expression {
    //   value: depth(SitesHierarchySimplified:^hierarchy) >= 1
    // }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_dnlistens), SitesHierarchySimplified:^hierarchy) > 0

    }
    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row selectedFlat #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      labelStyle: nodeOnly
    //showTotal: true
    }

    column #column_current_counts {
      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
      }

    }

    column #column_current_NPS {
      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
       // target: parseReal(SitesHierarchy:NPSTarget)
        navigateTo: page_DNListensResponses
       //view: comparativeStatisticView
      }
    }

    column #column_NPSGoal {

      label: "NPS® Goal"

      format: noDecimalNumber

      cell {
        value: parseReal(SitesHierarchySimplified:NPSTarget)
        //value: average(numeric(Goals_CustomTable:nps_target))
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_NPS_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_NPS
        other: column_NPSGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column cut #column_Promoters {

      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_DNListensResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_DNListensResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }
    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

      }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs_2 {
    label: "Location KPIs (hidden)"
    size: large
    hide: true
  //ignoreFilters: reportingPeriodFilter
    removeEmptyRows: true
    description: "### For Travel Hospitality, our NPS target is 61

Note: Overall Satisfaction measure included in survey starting April 27, 2023"


    select #Locations_Timeframe_Selector {
      label: "Select Timeframe for Trends"

      options: @valueSet_date_ranges_1.items
    } // end selector
    row cut #row_2 {
      value: :LocationName
      total: "none"
    }

    column {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber

      }

    }

    column {

      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        target: @reportConfig.nps_travel_target
        navigateTo: page_DNListensResponses
        view: comparativeStatisticView
      }
    }

    column cut {

      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_DNListensResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column {
      label: "NPS® Trends"
      filter expression {
        value: @Locations_Timeframe_Selector.selected.selectFilter
      }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Locations_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

    column #column_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_DNListensResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }
    column #column_OSAT_Trends {

      filter expression {
        value: @Locations_Timeframe_Selector.selected.selectFilter
      }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Locations_Timeframe_Selector.selected.selectBreakdownBy
        }

      }

      label: "Satisfaction Trends"
    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }
  } // end widget
  // widget keyDrivers #keyDriversWidget_OSAT_Travel {
  //   label: "What Drives Guest Satisfaction?"
  //   algorithm: regression
  //   dependentVariable: @reportConfig.osat_qid
  //   independentVariables: surveyDataset:SAT_DRIVERS.quality, surveyDataset:SAT_DRIVERS.value, surveyDataset:SAT_DRIVERS.variety, surveyDataset:SAT_DRIVERS.speed, surveyDataset:SAT_DRIVERS.staff
  //   satisfactionLimit: 85
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   quadrantColors: @reportConfig.kda_quadrantColors
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_regression
  //     info: @reportConfig.kda_infobox_info_regression
  //   }
  //   description: "This analysis looks for patterns in the data to determine how guest ratings on certain experiences influence their overall satisfaction with their visit. This shows us where to target improvement initiatives."
  //   importanceLimit: 0.2
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_OSAT_Travel
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments with Text Analytics**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  }
  widget comments #commentsWidget_Dining {
    label: "Comments with Text Analytics sentiment and categories"
    size: large
    table: textAnalyticsDataset_Dining.overallScore:
    sortOrder: descending
    sortColumn: responseColumn

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000
    navigateTo: page_Indiv_Survey_Response_TA

    infobox #infobox {
      label: "Information"
      info: "This widget shows all verbatim comments, and the comment's overall sentiment or other contextual variables related to the comment. 
- Overall sentiment is measured for all the text in a comment field rather than parts of it.
- Overall sentiment ranges from -5 to 5. 0 is neutral or mixed. 
- Tags under each comment represent the topic categories associated with this comment. Tags are color-coded red for negative, yellow for neutral/mixed and green for positive. 
- Columns are filterable.
- Clicking anywhere on a comment will bring you to the Response-level results."
    }


    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: large
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: large
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
    }

    group question #questionGroup {
      label: "All Comments"
      comment: textAnalyticsDataset_Dining.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Dining.overallScore:text != ""
      }
    }
    column response #responseColumn {
      sortBy: footer
      //header: "Claim #" + surveyDataset:ClaimNbr
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta

      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "Comment Field"
      value: textAnalyticsDataset_Dining.overallScore:variable
      enableColumnFilter: true
      width: 150px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #StoreName {
      label: "Store / Restaurant"
      value: surveyDataset_TA:STORE_INFO
      enableColumnFilter: true
      //value: surveyDataset_TA:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Dining:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Dining:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 125px
    }

    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    column metric #metricColumn_NPS {
      label: "NPS"
      value: score(@reportConfig.nps_qid_ta)
      enableColumnFilter: true
      //filterable: true
      width: 125px
      align: center
      view: colorcoding
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_OSAT {
      label: "SAT"
      value: score(@reportConfig.osat_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }


    description: "**Note: To filter on Overall Sentiment, enter 3 for Positive, 2 for Neutral, 1 for Negative**
    **Note: To filter on NPS Segment, enter 3 for Promoters, 2 for Passives, 1 for Detractors**"


  } // end widget
  widget chart #TopTopics_chartWidget {

  //  label: @TANumTopics_Selector.selectedLabel + " " + @TACategoryLevels_Selector.selectedLabel + " by Volume"
    label: "Top 10 Text Analytics Topics by Volume"

    size: large
    animation: false
    gridLines: false
    legend: bottomCenter
    layout: "horizontal"
    palette: palettePosNegNueReverse

    hide: false

    filter expression {
      //value: depth(textAnalyticsDataset_Dining.model:^parent) = @TACategoryLevels_Selector.selected
      value: depth(textAnalyticsDataset_Dining.model:^parent) = 1
    }

    series #volume1 {
      label: "Mentions"
      value: textAnalyticsDataset_Dining:categoryCountTASet1()
      format: noDecimalNumber
      //navigateFilter: some(textAnalyticsDataset_Dining.categoryScore:, true, textAnalyticsDataset_Dining.categoryScore:)
      //navigateTo: dd_CategoryResultsByThemeComments
      navigateTo: dd_SentimentComments_Dining

      breakdownBy cut {
        value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      }
      percent: false
      chart bar {
        mode: stacked
        maxBarSize: 65
      }
    }
    category selectedFlat {
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
     // takeTop: @TANumTopics_Selector.selected
      takeTop: 10
      sortBy: "volume1"
      sortOrder: descending
    }


    axis secondary {
      label: "Category Sentiment"
      hide: true
    }

    axis category #categoryAxis {

      textSize: 150
      orientation: "-45"
    }
    axis primary {
      format: noDecimalNumber
    }
    navigateTo: "page_Parks_Overview"
  } // end widget
  // widget headline #headlineWidget_8 {
  //   label: "Text Analytics Sentiment Trends"
  //   size: large
  //   cardBackground: @reportConfig.selector_CardBackgroundColor


  //   select #TA_Timeframe_Selector_Dining {
  //     label: "Select a Timeframe"
  //     options: @valueSet_date_ranges.items

  //   } // end selector
  //   tile markdown #markdownTile {
  //     value: "### The section displays sentiment trends."
  //   }

  // } // end widget
  widget chart #SentimentTrends_chartWidget {
    label: "Text Analytics Sentiment Components Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    size: large
    animation: true
    gridLines: horizontal
    legend: bottomCenter
    removeEmptyCategories: true
    hide: true
    //navigateTo: dd_SentimentComments
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Timeframe_SelectorTA1.selected.selectFilter
    // }

    infobox #infobox {
      label: "Information"
      info: "This widget shows the % distribution of overall sentiment over time. Time period break (first drop-down menu) and sentiment group base (second drop-down menu) may be selected. The distribution of the sentiment group is based on either respondents or comments for (All, positive, neutral/mixed, or negative). 
- Overall sentiment is measured for all the text in a comment field rather than parts of it. 
- Hover over the dots for more info.
- Clicking on a bar or dot will take you to the category results for that time period."
    }

    series #series_primary {
      chart bar {
        mode: "stacked100Percent"
        dataLabel: percentThenValue
        barSize: 75
        maxBarSize: 75
      }
      value: textAnalyticsDataset_Dining:overallResponseBaseTASet1()
      label: "% distribution of respondents by sentiment group"
      format: noDecimalNumber
     // format: @metric_selector.selected.cellFormat
      palette: paletteNegNeuPos
      navigateTo: dd_SentimentComments_Dining

      breakdownBy cut #cutBreakdownby {
        value: textAnalyticsDataset_Dining:responseSentimentGroup()
      }
    }

    series #series_secondary {
      value: textAnalyticsDataset_Dining:overallAverageTASet1()
      format: oneDecimalNumber
      label: "Average Sentiment"
      isSecondary: true
      chart line {
        lineWidth: 3
        dotSize: 7
        dotColorFormat: taSentimentColorDefaultFormatter
        connectNulls: true
        showDotValue: true
      }
      palette: palettePosNegNueReverse
    }


    category date #cutByDate {
      value: @reportConfig.intvdate_ta
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

    }

    chartMargin {
      top: 20
    }
    axis primary {
      label: "%"
      format: percentNoDecimal
      minValue: 0
      maxValue: 100
    }
    axis category {
      orientation: -45
      textSize: 75
    }
    axis secondary #secondaryAxis {
      label: "Sentiment (-5 to 5)"
      minValue: -5
      maxValue: 5
      format: noDecimalNumber
    }
    base {
      value: textAnalyticsDataset_Dining:overallResponseBaseTASet1()
      format: baseNumberFormatter
    }
    removeEmptySeries: true
  } // end widget
  widget headline #CatsAndSentiment_headlineWidget {
    label: "Text Analytics Categories & Sentiment Analysis"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #HierView_Selector {
      label: "Select a View"
      options: @valueSet_hierarchy_views.items

    } // end selector
    tile markdown #markdownTile {
      value: "###"
    }

  } // end widget
  widget dataGrid #CatsAndSentiment_HierView {
    label: "Text Analytics Categories & Sentiment - Hierarchical View"
    size: "large"

    hide: @HierView_Selector.selected != 1

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedHierarchy #comparisonRow {
      sortBy: "/percentTotalComments"
      sortOrder: descending
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:percentageOfCommentsTASet1()
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Dining:categoryCountTASet1()
        format: noDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

        }
        format: oneDecimalNumber

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Dining:categoryCount()
        extraValue: textAnalyticsDataset_Dining:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
  widget dataGrid #CatsAndSentiment_FlatView {
    label: "Text Analytics Categories & Sentiment - Flat view"
    size: "large"
    //navigateTo: dd_CategoryResultsByThemeComments

    hide: @HierView_Selector.selected != 2

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector


    row selectedFlat #comparisonRow {
      sortOrder: descending
      sortBy: "/percentTotalComments"
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:percentageOfCommentsTASet1()
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Dining:categoryCountTASet1()
        format: noDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Microcharts_Timeframe_Selector.selected.selectFilter
      // }
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()

        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

        }
        format: oneDecimalNumber

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Dining:categoryCount()
        extraValue: textAnalyticsDataset_Dining:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }

    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }
  } // end widget
  widget markdown #markdownWidget_PerformanceTrends {
    markdown: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    size: large
  }
  widget dataGrid #dataGridWidget_SatDrivers {
    label: "Satisfaction Drivers"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_DRIVERS$field
      total: none

    }
    column #column_current_counts {
      value: count(:SAT_DRIVERS$value)
      label: "Number of Responses"
      cell {
        value: count(:SAT_DRIVERS$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

    description: "Note: Variety and Value measures included in survey starting April 27, 2023.  Quality, Speed of Service, and Friendliness of Staff were included in the survey starting February 6, 2023.

Note: 'N/A' responses have been filtered out of the results below."
  } //end widget
  widget dataGrid #dataGridWidget_Sat_TimeOfDay {
    label: "Satisfaction By Time of Day"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    // sort rows {
    //   sortBy: "/Satisfaction"
    //   sortOrder: descending
    // }

    row cut {
      value: surveyDataset:TIME_OF_VISIT
      total: none

    }
    column #column_current_counts {
      value: count(surveyDataset:TIME_OF_VISIT)
      label: "Number of Responses"
      cell {
        value: count(surveyDataset:TIME_OF_VISIT)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }


    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023"
  } //end widget
  // widget chart #dataGridWidget_Sat_TimeOfVisit {
  //   label: "Satisfaction By Time of Visit" + " - " + @Travel_Timeframe_Selector.selectedLabel
  //   // label: @kpiselect.selected.kpiLabel + " Trends"   
  //   palette: multicolors1_palette
  //  // ignoreFilters: reportingPeriodFilter

  //   // select #TimeofDay_Timeframe_Selector {
  //   //   label: "Select Timeframe"

  //   //   options: @valueSet_date_ranges_1.items

  //   // } // end selector
  //   size: halfwidth

  //   legend: bottomCenter
  //   chartMargin {
  //     top: 20
  //     bottom: 75
  //     right: 25
  //   }

  //   series #series {
  //     chart line {
  //       showDotValue: false

  //     }

  //     value: top1percent(@reportConfig.osat_qid)
  //     format: oneDecimalPercent

  //     isSecondary: false
  //     breakdownBy cut {
  //       value: surveyDataset:TIME_OF_VISIT

  //     }
  //   }

  //   category date #dateCategory {
  //     value: @reportConfig.intvdate
  //     breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
  //     label: "Interview date"
  //     //format: dateDefaultFormatter
  //   }


  //   axis category #categoryAxis {
  //     orientation: "-45"
  //     format: noDecimalPercent

  //   }
  //   axis primary #primaryAxis {
  //        //  format: metricsItemMetricDefaultFormatter
  //     format: noDecimalPercent
  //     label: "% Very Satisfied"
  //     minValue: 50
  //     maxValue: 100
  //   }
  //   axis secondary #secondaryAxis {
  //     hide: true
  //     label: "% Response"
  //     format: noDecimalPercent
  //     minValue: 0
  //     maxValue: 100
  //   }


  //   base #base {
  //     value: count(@reportConfig.osat_qid)
  //     format: baseNumberFormatter
  //   }
  //   removeEmptyCategories: true
  //   removeEmptySeries: true
  // } // end widget
} // end page
page #page_Lodging_Overview {
  label: "Parks & Resorts - Lodging"

  access rules {
    rule claim {
      name: "UserSegment"
      value: "All", "Lodging", "Parks"
      //value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_LodgingSurvey()
    label: "Lodging survey Only"
  }


  filter expression #NPSAnswered2 {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  filter expression {
    value: surveyDataset:filterMeasure_ExcludeAustraliaLocations()
    label: "Exclude Australia locations"
  }

  widget headline #headlineWidget_Lodging_Overview {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Parks & Resorts - Lodging 
### This dashboard compiles lodging survey data collected  via emails sent directly to guests within 1 day post visit. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatim comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a location. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }

    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }

    tile button #buttonTile {
      value: "Click here to see information about guest demographics"
      navigateTo: "page_Demos"
      navigateOptions: "same_tab"

      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
    }
    label: "Voice of Guest Dashboard"
  }
  widget kpi #kpiWidget_Overall_NPS {
    label: "Overall Subsidiary NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
     // target: @reportConfig.nps_lodging_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all lodging locations with Parks & Resorts.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Overall Subsidiary OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_lodging_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all lodging locations with Parks & Resorts.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Parks & Resorts location(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small


    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Parks & Resorts location(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }



  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  }

  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_LodgingSurvey()
      type: primary


      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_LodgingSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_LodgingSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
    }
  }
  widget headline #headlineWidget_totalOpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :PROBLEM
    }
    palette: redtogreen2ptscale

    navigateTo: "page_Parks_Overview"
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  }
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Lodging_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @NPS_Timeframe_Selector2.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector2 {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent

        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal
      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter

    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @OSAT_Timeframe_Selector2.selected.selectFilter
    // }

    // select #OSAT_Timeframe_Selector2 {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "This view displays a breakdown of the performance of all locations on our key performance indicators. This provides insight on how locations perform in a relative context.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_lodging), SitesHierarchySimplified:^hierarchy) > 0

    }

    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_current_counts {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        navigateTo: page_LodgingResponses

      }

    }

    column #column_current_NPS {

      label: "NPS®"

      // scope reportingPeriod {
      //   period: Current
      // }
      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        navigateTo: page_LodgingResponses
       // view: comparativeStatisticView
      }
    }

    column cut #column_Promoters {
      //value: recode(@reportConfig.nps_qid, @NPScats)
      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_LodgingResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Lodging_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_current_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_LodgingResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }

    column #column_OSATGoal {

      label: "OSAT Goal"

      format: noDecimalNumber

      cell {

        value: parseReal(SitesHierarchySimplified:OSATTarget)
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_OSAT_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_OSAT
        other: column_OSATGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Lodging_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        }

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget headline #headlineWidget_KDAs_Location {
    label: "Key Driver Analysis By Location"
    size: large

    tile markdown #markdown1 {
      value: "### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

### The data below show the relationships at high levels as well as at functional levels."

//### **Please note:** These analyses require a minimum of 100 records to run; if less than 100 records are available, the report will generate an error message. If you see the message 'The accuracy of the model shown falls below the criteria specified. Please exercise caution in the use of these data.' this means that the R-squared value of the model falls below 0.5."

    }

    select #Lodging_Locations_Selector {
      label: "Select a Lodging Location"

      options: @valueSet_lodging_locations.items

    } // end selector
  }
//   widget markdown #markdownWidget_3 {
//     markdown: "## **Key Driver Analysis**

// ### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

// ### The data below show the relationships at high levels as well as at functional levels. "
//     size: large
//   }

  // widget keyDrivers #keyDriversWidget_NPS_Lodging_Overall {
  //   label: "What Drives Likelihood to Recommend for Lodging Overall?"

  // //attributes removed for this KDA: none
  // //this kda applies to lodging as a whole

  //   hide: @Lodging_Locations_Selector.selected != "Lodging"
  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

  //   minimumSampleSize: @reportConfig.KDAMinimumSampleSize
  //   algorithm: correlation
  //   satisfactionLimit: 80
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: @reportConfig.kda_descriptionText
  //   importanceLimit: 0.5
  //   dependentVariable: surveyDataset:NPS
  //   independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.concierge, surveyDataset:SAT_EXPERIENCES.otheramenities, surveyDataset:SAT_EXPERIENCES.spa, surveyDataset:SAT_EXPERIENCES.shops

  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_NPS_Lodging_Overall

  widget keyDrivers #keyDriversWidget_NPS_Lodging1 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

  //attributes removed for this KDA: breakfast
  //this kda applies to following locations:
    //474A	The Lodge at Tenaya 
    //474B	The Cottages at Tenaya
    //474C	The Explorer Cabins at Tenaya  

    hide: @Lodging_Locations_Selector.selected != "474A" AND @Lodging_Locations_Selector.selected != "474B" AND @Lodging_Locations_Selector.selected != "474C"
    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.concierge, surveyDataset:SAT_EXPERIENCES.otheramenities, surveyDataset:SAT_EXPERIENCES.spa, surveyDataset:SAT_EXPERIENCES.shops

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging1
  widget keyDrivers #keyDriversWidget_NPS_Lodging2 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, spa, other amenities
   //this kda applies to following locations:
    //59841	Peaks of Otter
    //59989A	John Muir Lodge - Kings Canyon National Park
    //59989B	Grant Grove Cabins - Kings Canyon National Park
    //63108	Yavapai Lodge - Grand Canyon National Park
    //63275	Trailer Village RV Park - Grand Canyon National Park

    hide: @Lodging_Locations_Selector.selected != "59841" AND @Lodging_Locations_Selector.selected != "59989A" AND @Lodging_Locations_Selector.selected != "59989B" AND @Lodging_Locations_Selector.selected != "63108" AND @Lodging_Locations_Selector.selected != "63275"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.shops

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging2
  widget keyDrivers #keyDriversWidget_NPS_Lodging3 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, spa
   //this kda applies to following locations:
    //22005A	The Lodge at Geneva on the Lake
    //22005B	The Cottages at Geneva on the Lake
    //58866	Big Meadows Lodge - Shenandoah
    //58867	Skyland Resort - Shenandoah

    hide: @Lodging_Locations_Selector.selected != "22005A" AND @Lodging_Locations_Selector.selected != "22005B" AND @Lodging_Locations_Selector.selected != "58866" AND @Lodging_Locations_Selector.selected != "58867"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.shops, surveyDataset:SAT_EXPERIENCES.otheramenities

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging3
  widget keyDrivers #keyDriversWidget_NPS_Lodging4 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, spa, bars, other amenities
   //this kda applies to following locations:
    //404	Wuksachi Lodge - Sequoia National Park   
    //58148	Kalaloch Lodge
    //59988	Cedar Grove Lodge - Kings Canyon National Park

    hide: @Lodging_Locations_Selector.selected != "404" AND @Lodging_Locations_Selector.selected != "58148" AND @Lodging_Locations_Selector.selected != "59988"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.shops

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging4
  widget keyDrivers #keyDriversWidget_NPS_Lodging5 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, bars, other amenities
   //this kda applies to following locations:
    //139	The Gideon Putnam

    hide: @Lodging_Locations_Selector.selected != "139"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.shops, surveyDataset:SAT_EXPERIENCES.spa

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging5
  widget keyDrivers #keyDriversWidget_NPS_Lodging6 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: concierge, restaurants, bars, shops, spa
   //this kda applies to following locations:
    //28577	Gray Wolf Inn & Suites
    //28578	Yellowstone Park Hotel


    hide: @Lodging_Locations_Selector.selected != "28577" AND @Lodging_Locations_Selector.selected != "28578"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.breakfast, surveyDataset:SAT_EXPERIENCES.otheramenities

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging6
  widget keyDrivers #keyDriversWidget_NPS_Lodging7 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, restaurants, bars, shops, spa
   //this kda applies to following locations:
    //59396	The Explorer Cabins at Yellowstone

    hide: @Lodging_Locations_Selector.selected != "59396"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.otheramenities

    warningText: @reportConfig.kda_warningText
    //rSquaredLimit: 0.5
  } // end widget keyDriversWidget_NPS_Lodging7
  widget headline #headlineWidget_KDAs_Location_Addtl {

    label: "Additional Key Driver Analyses for " + @Lodging_Locations_Selector.selectedLabel + ""
    size: large

    select #lodging_addl_keydrivers_selector {
      label: "Select an Additional Key Driver Analysis"
      options: item {
        label: "Select to see other Key Driver Analyses"
        value: 0
      },
      item {
        label: "What Drives Satisfaction with Lodging?"
        value: 1
      },
      item {
        label: "How Do Room Features Impact Lodging Satisfaction?"
        value: 2
      },
      item {
        label: "What Drives Restaurant Satisfaction?"
        value: 3
      },
      item {
        label: "What Drives Bar Satisfaction?"
        value: 4
      }

    }

    tile markdown #markdownTile_2 {
      value: "### There are several analytic views that provide us with strategic direction on what areas to promote as well as those areas that we should consider fixing . To view these, please select  an analysis from the dropdown above."
    }

  }

  // widget keyDrivers #keyDriversWidget_SAT_Lodging_Overall {
  //   label: "What Drives Satisfaction with Lodging Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 1 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

  //   minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    // algorithm: regression
    //// algorithm: correlation

  //   satisfactionLimit: 85
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
  //   importanceLimit: 0.15
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
  //   independentVariables: surveyDataset:DRILL_LODGING.accuracy, surveyDataset:DRILL_LODGING.arrival, surveyDataset:DRILL_LODGING.avail, surveyDataset:DRILL_LODGING.cleanliness, surveyDataset:DRILL_LODGING.staff, surveyDataset:DRILL_LODGING.departure, surveyDataset:DRILL_LODGING.service
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Lodging_Overall

  widget keyDrivers #keyDriversWidget_SAT_Lodging {
    label: "What Drives Satisfaction with Lodging at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 1

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
    independentVariables: surveyDataset:DRILL_LODGING.accuracy, surveyDataset:DRILL_LODGING.arrival, surveyDataset:DRILL_LODGING.avail, surveyDataset:DRILL_LODGING.cleanliness, surveyDataset:DRILL_LODGING.staff, surveyDataset:DRILL_LODGING.departure, surveyDataset:DRILL_LODGING.service
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Lodging
  // widget keyDrivers #keyDriversWidget_SAT_Room_Overall {
  //   label: "How Do Room Features Impact Lodging Satisfaction Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 2 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

    // algorithm: regression
    //// algorithm: correlation
  //   satisfactionLimit: 85
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how room features, experiences and characteristics influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
  //   importanceLimit: 0.10
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
  //   independentVariables: surveyDataset:DRILL_ROOM.ac, surveyDataset:DRILL_ROOM.bathamenities, surveyDataset:DRILL_ROOM.bathclean, surveyDataset:DRILL_ROOM.bathfeatures, surveyDataset:DRILL_ROOM.bed, surveyDataset:DRILL_ROOM.cleanliness, surveyDataset:DRILL_ROOM.furnishings, surveyDataset:DRILL_ROOM.quiet, surveyDataset:DRILL_ROOM.smell, surveyDataset:DRILL_ROOM.wifi
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Room_Overall

  widget keyDrivers #keyDriversWidget_SAT_Room {
    label: "How Do Room Features Impact Lodging Satisfaction at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 2

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how room features, experiences and characteristics influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
    independentVariables: surveyDataset:DRILL_ROOM.ac, surveyDataset:DRILL_ROOM.bathamenities, surveyDataset:DRILL_ROOM.bathclean, surveyDataset:DRILL_ROOM.bathfeatures, surveyDataset:DRILL_ROOM.bed, surveyDataset:DRILL_ROOM.cleanliness, surveyDataset:DRILL_ROOM.furnishings, surveyDataset:DRILL_ROOM.quiet, surveyDataset:DRILL_ROOM.smell, surveyDataset:DRILL_ROOM.wifi
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Room
  // widget keyDrivers #keyDriversWidget_SAT_Restaurants_Overall {
  //   label: "What Drives Restaurant Satisfaction Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 3 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

  //   select #catfilter {
  //     label: "Filter by Meal Rated"
  //     mode: multi

  //     options: @categorySet_meal_rated.items
  //   }
  //   filter expression {
  //     value: selected(:MEAL_RATED, @catfilter.selected)
  //   }

    // algorithm: regression
    //// algorithm: correlation
  //   satisfactionLimit: 80
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
  //   importanceLimit: 0.15
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.restaurants
  //   independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Restaurants_Overall

  widget keyDrivers #keyDriversWidget_SAT_Restaurants {
    label: "What Drives Restaurant Satisfaction at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 3

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    select #catfilter {
      label: "Filter by Meal Rated"
      mode: multi

      options: @categorySet_meal_rated.items
    }
    filter expression {
      value: selected(:MEAL_RATED, @catfilter.selected)
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation

      size: large
    }
    description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_EXPERIENCES.restaurants
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Restaurants
  // widget keyDrivers #keyDriversWidget_SAT_Bars_Overall {
  //   label: "What Drives Bar Satisfaction Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 4 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }
  //   minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    // algorithm: regression
    //// algorithm: correlation
  //   satisfactionLimit: 86
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the bar influence their overall bar satisfaction. This shows us where to target improvement in our bar processes and experiences."
  //   importanceLimit: 0.10
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.bars
  //   independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Bars_Overall

  widget keyDrivers #keyDriversWidget_SAT_Bars {
    label: "What Drives Bar Satisfaction at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 4

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 86
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the bar influence their overall bar satisfaction. This shows us where to target improvement in our bar processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT_EXPERIENCES.bars
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Bars
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments with Text Analytics**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  }



   //begin TA Lodging
  widget comments #commentsWidget1 {
    label: "Comments with Text Analytics sentiment and categories"
    size: large
    table: textAnalyticsDataset_Lodging.overallScore:
    sortOrder: descending
    sortColumn: responseColumn

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response_TA

    infobox #infobox {
      label: "Information"
      info: "This widget shows all verbatim comments, and the comment's overall sentiment or other contextual variables related to the comment. 
- Overall sentiment is measured for all the text in a comment field rather than parts of it.
- Overall sentiment ranges from -5 to 5. 0 is neutral or mixed. 
- Tags under each comment represent the topic categories associated with this comment. Tags are color-coded red for negative, yellow for neutral/mixed and green for positive. 
- Columns are filterable.
- Clicking anywhere on a comment will bring you to the Response-level results."
    }


    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
      fontSize: medium
    }

    group question #questionGroup {
      label: "All Comments"
      comment: textAnalyticsDataset_Lodging.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Lodging.overallScore:text != ""
      }
    }
    column response #responseColumn {
      sortBy: footer
      //header: "Claim #" + surveyDataset:ClaimNbr
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta

      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "Comment Field"
      value: textAnalyticsDataset_Lodging.overallScore:variable
      enableColumnFilter: true
      width: 150px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Lodging:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Lodging:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 125px
    }

    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    column metric #metricColumn_NPS {
      label: "NPS"
      value: score(@reportConfig.nps_qid_ta)
      enableColumnFilter: true
      //filterable: true
      width: 125px
      align: center
      view: colorcoding
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_OSAT {
      label: "SAT"
      value: score(@reportConfig.osat_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }


    description: "**Note: To filter on Overall Sentiment, enter 3 for Positive, 2 for Neutral, 1 for Negative**
    **Note: To filter on NPS Segment, enter 3 for Promoters, 2 for Passives, 1 for Detractors**"


  } // end widget
  widget chart #TopTopics_chartWidget {

  //  label: @TANumTopics_Selector.selectedLabel + " " + @TACategoryLevels_Selector.selectedLabel + " by Volume"
    label: "Top 10 Text Analytics Topics by Volume"

    size: large
    animation: false
    gridLines: false
    legend: bottomCenter
    layout: "horizontal"
    palette: palettePosNegNueReverse

    hide: false

    filter expression {
      //value: depth(textAnalyticsDataset_Lodging.model:^parent) = @TACategoryLevels_Selector.selected
      value: depth(textAnalyticsDataset_Lodging.model:^parent) = 2
    }

    series #volume1 {
      label: "Mentions"
      value: textAnalyticsDataset_Lodging:categoryCountTASet1()
      format: noDecimalNumber
      //navigateFilter: some(textAnalyticsDataset_Lodging.categoryScore:, true, textAnalyticsDataset_Lodging.categoryScore:)
      //navigateTo: dd_CategoryResultsByThemeComments
      navigateTo: dd_SentimentComments_Lodging

      breakdownBy cut {
        value: textAnalyticsDataset_Lodging.categoryScore:categorySentimentGroup
      }
      percent: false
      chart bar {
        mode: stacked
        maxBarSize: 65
      }
    }
    category selectedFlat {
      reportingHierarchy: textAnalyticsDataset_Lodging:categoryHierarchy_Lodging
     // takeTop: @TANumTopics_Selector.selected
      takeTop: 10
      sortBy: "volume1"
      sortOrder: descending
    }


    axis secondary {
      label: "Category Sentiment"
      hide: true
    }

    axis category #categoryAxis {

      textSize: 100
      orientation: "-45"
    }
    axis primary {
      format: noDecimalNumber
    }
    navigateTo: "page_Parks_Overview"
  } // end widget
  // widget headline #SentimentTrends_headlineWidget {
  //   label: "Text Analytics Sentiment Trends"
  //   size: large
  //   cardBackground: @reportConfig.selector_CardBackgroundColor


  //   select #Timeframe_SelectorTA1 {
  //     label: "Select a Timeframe"
  //     options: @valueSet_date_ranges.items

  //   } // end selector
  //   tile markdown #markdownTile {
  //     value: "### The section displays sentiment trends."
  //   }

  // } // end widget
  widget chart #SentimentTrends_chartWidget {
    label: "Text Analytics Sentiment Components Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
    size: large
    animation: true
    gridLines: horizontal
    legend: bottomCenter
    removeEmptyCategories: true
    //navigateTo: dd_SentimentComments
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Timeframe_SelectorTA1.selected.selectFilter
    // }

    infobox #infobox {
      label: "Information"
      info: "This widget shows the % distribution of overall sentiment over time. Time period break (first drop-down menu) and sentiment group base (second drop-down menu) may be selected. The distribution of the sentiment group is based on either respondents or comments for (All, positive, neutral/mixed, or negative). 
- Overall sentiment is measured for all the text in a comment field rather than parts of it. 
- Hover over the dots for more info.
- Clicking on a bar or dot will take you to the category results for that time period."
    }

    series #series_primary {
      chart bar {
        mode: "stacked100Percent"
        dataLabel: percentThenValue
        barSize: 75
        maxBarSize: 75
      }
      value: textAnalyticsDataset_Lodging:overallResponseBaseTASet1()
      label: "% distribution of respondents by sentiment group"
      format: noDecimalNumber
     // format: @metric_selector.selected.cellFormat
      palette: paletteNegNeuPos
      navigateTo: dd_SentimentComments_Lodging

      breakdownBy cut #cutBreakdownby {
        value: textAnalyticsDataset_Lodging:responseSentimentGroup()
      }
    }

    series #series_secondary {
      value: textAnalyticsDataset_Lodging:overallAverageTASet1()
      format: oneDecimalNumber
      label: "Average Sentiment"
      isSecondary: true
      chart line {
        lineWidth: 3
        dotSize: 7
        dotColorFormat: taSentimentColorDefaultFormatter
        connectNulls: true
        showDotValue: true
      }
      palette: palettePosNegNueReverse
    }


    category date #cutByDate {
      value: @reportConfig.intvdate_ta
      breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    chartMargin {
      top: 20
    }
    axis primary {
      label: "%"
      format: percentNoDecimal
      minValue: 0
      maxValue: 100
    }
    axis category {
      orientation: -45
      textSize: 75
    }
    axis secondary #secondaryAxis {
      label: "Sentiment (-5 to 5)"
      minValue: -5
      maxValue: 5
      format: noDecimalNumber
    }
    base {
      value: textAnalyticsDataset_Lodging:overallResponseBaseTASet1()
      format: baseNumberFormatter
    }
    removeEmptySeries: true
  } // end widget
  widget headline #CatsAndSentiment_headlineWidget {
    label: "Text Analytics Categories & Sentiment Analysis"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #HierView_Selector {
      label: "Select a View"
      options: @valueSet_hierarchy_views.items

    } // end selector
    tile markdown #markdownTile {
      value: "###"
    }

  } // end widget
  widget dataGrid #CatsAndSentiment_HierView {
    label: "Text Analytics Categories & Sentiment - Hierarchical View"
    size: "large"

    hide: @HierView_Selector.selected != 1

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedHierarchy #comparisonRow {
      sortBy: "/percentTotalComments"
      sortOrder: descending
      reportingHierarchy: textAnalyticsDataset_Lodging:categoryHierarchy_Lodging
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Lodging:percentageOfCommentsTASet1()
        format: percentNoDecimal
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Lodging
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Lodging:categoryCountTASet1()
        format: noDecimalNumber

        navigateTo: dd_SentimentComments_Lodging
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Lodging:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber

        navigateTo: dd_SentimentComments_Lodging
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
      filter expression {
        value: @Lodging_Timeframe_Selector.selected.selectFilter
      }
      cell microchart #cell {
        value: textAnalyticsDataset_Lodging:categoryAverageTASet1()
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
          align: true
          //start: "-4 quarter"

        }
        format: oneDecimalNumber

      }

    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Lodging.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Lodging:categoryCount()
        extraValue: textAnalyticsDataset_Lodging:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal

        navigateTo: dd_SentimentComments_Lodging
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
  widget dataGrid #CatsAndSentiment_FlatView1 {
    label: "Text Analytics Categories & Sentiment - Flat view"
    size: "large"


    hide: @HierView_Selector.selected != 2

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedFlat #comparisonRow {
      sortOrder: descending
      sortBy: "/percentTotalComments"
      reportingHierarchy: textAnalyticsDataset_Lodging:categoryHierarchy_Lodging
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Lodging:percentageOfCommentsTASet1()
        format: percentNoDecimal
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Lodging
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Lodging:categoryCountTASet1()
        format: noDecimalNumber
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Lodging
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Lodging:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Lodging
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends"

      cell microchart #cell {
        value: textAnalyticsDataset_Lodging:categoryAverageTASet1()

        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
          align: true
          //start: "-4 quarter"
        }
        format: oneDecimalNumber

      }

    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Lodging.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Lodging:categoryCount()
        extraValue: textAnalyticsDataset_Lodging:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal

        navigateTo: dd_SentimentComments_Lodging
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
  widget headline #headlineWidget_15 {

    label: ""
    size: large
    hide: true
    tile markdown #markdownTile_2 {
      value: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    }

  }
  widget chart #chartWidget_NPS_Trends_Lines {
    label: "NPS® Trends"
    hide: true
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
    // ignoreFilters: reportingPeriod

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series1 {
      chart line {
        showDotValue: true

      }

      value: nps(@reportConfig.nps_qid) * 100
      format: noDecimalNumber
      label: "NPS®"

    }

    series #series2 {
      chart line {
        showDotValue: false

      }

      percentOver: series
      value: count(@reportConfig.nps_qid)
      format: oneDecimalPercent

      isSecondary: true
      breakdownBy cut {
        value: :NPSVal

      }
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 75
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Lines {
    label: "Overall Satisfaction (Top Box) Trend"
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
    hide: true
    // ignoreFilters: reportingPeriod
    // hide: false

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series1 {
      chart line {
        showDotValue: true

      }

      value: top1percent(@reportConfig.osat_qid)
      format: oneDecimalPercent
      label: "Overall Satisfaction"

    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: oneDecimalPercent
      label: "Top Box % (5's)"
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "% Response"
      format: noDecimalPercent
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      right: 20
      bottom: 75
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
  } // end widget
  widget markdown #markdownWidget_PerformanceTrends {
    markdown: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    size: large
  }
  widget dataGrid #dataGridWidget_ExperiencesSat {
    label: "Satisfaction with Experiences"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_EXPERIENCES$field
      total: none

    }
    column #column_current_counts {

      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:SAT_EXPERIENCES$value)

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell #undefined {
        format: noDecimalPercent
        value: top1percent(:SAT_EXPERIENCES$value)
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_EXPERIENCES$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_LodgingSat {
    label: "Lodging Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_LODGING$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_LODGING$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_LODGING$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RoomSat {
    label: "Room Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_ROOM$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_ROOM$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_ROOM$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RestaurantSat {
    label: "Restaurant Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    select #catfilter {
      label: "Filter by Meal Rated"
      mode: multi

      options: @categorySet_meal_rated.items
    }
    filter expression {
      value: selected(:MEAL_RATED, @catfilter.selected)
    }

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_RESTAURANT$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_RESTAURANT$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_RESTAURANT$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RVParkSat {
    label: "RV Park Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }


    row cut {
      value: :DRILL_TRAILER_PARK$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_TRAILER_PARK$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_TRAILER_PARK$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_TRAILER_PARK$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }


  } //end widget
  widget headline #headlineWidget_LocationKPISummaries {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "# **Location-Based KPI Summaries**
### This section looks at how specific locations track on our KPI's (and the trends)."
    }

  }
  widget dataGrid #dataGridWidget_LocationPerfTrends {
    label: "Location Performance Trends"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_Arrival {
      label: "Arrival (Top Box)"
      cell #cell {
        value: top1percent(:DRILL_LODGING.arrival)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        extraValue: count(:DRILL_LODGING.arrival)
        extraValueFormat: noDecimalNumber

        navigateTo: page_LodgingResponses
        navigateFilter: _isnotnull(:DRILL_LODGING.arrival)
      }

    }

    column #column_Arrival_Trends {
      label: "Arrival Sat Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
      cell microchart #cell {
        value: top1percent(:DRILL_LODGING.arrival)
        format: oneDecimalPercent
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }
      }

    }

    column #column_CleanRoom {
      label: "Clean Room (Top Box)"
      cell #cell {
        value: top1percent(:DRILL_ROOM.cleanliness)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        extraValue: count(:DRILL_ROOM.cleanliness)
        extraValueFormat: noDecimalNumber

        navigateTo: page_LodgingResponses
        navigateFilter: _isnotnull(:DRILL_ROOM.cleanliness)
      }

    }

    column #column_CleanRoom_Trends {
      label: "Clean Room Sat Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
      cell microchart #cell {
        value: top1percent(:DRILL_ROOM.cleanliness)
        format: oneDecimalPercent
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }
      }

    }

    column #column_CleanBathroom {
      label: "Clean Bathroom (Top Box)"
      cell #cell {
        value: top1percent(:DRILL_ROOM.bathclean)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        extraValue: count(:DRILL_ROOM.bathclean)
        extraValueFormat: noDecimalNumber

        navigateTo: page_LodgingResponses
        navigateFilter: _isnotnull(:DRILL_ROOM.bathclean)
      }

    }

    column #column_CleanBathroom_Trends {
      label: "Clean Bathroom Sat Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
      cell microchart #cell {
        value: top1percent(:DRILL_ROOM.bathclean)
        format: oneDecimalPercent
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }
      }

    }

    column #column_Restaurants {
      label: "Restaurants Sat (Top Box)"
      cell #cell {
        value: top1percent(:SAT_EXPERIENCES.restaurants)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        extraValue: count(:SAT_EXPERIENCES.restaurants)
        extraValueFormat: noDecimalNumber

        navigateTo: page_LodgingResponses
        navigateFilter: _isnotnull(:SAT_EXPERIENCES.restaurants)
      }

    }
    column #column_Restaurants_Trends {
      label: "Restaurants Sat Trends" + " - " + @Lodging_Timeframe_Selector.selectedLabel
      cell microchart #cell {
        value: top1percent(:SAT_EXPERIENCES.restaurants)
        format: oneDecimalPercent
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }
      }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: ""
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }
  } // end widget
  hide: false
  modal: false
} // end page
page #page_Tours_Overview {
  label: "Parks & Resorts - Tours"
  hide: false
  access rules {
    rule claim {
      name: "UserSegment"
      value: "All", "Tours", "Parks"
      //value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }

  layoutArea toolbar {
    filter multiselect #f_TourActivities {
      label: "Tour Activities"
      optionsFrom: :TourActivityName
    }
  }

  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_ToursSurvey()
    label: "Tours survey Only"
  }


  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }


  widget headline #headlineWidget_10 {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Tours 
### This dashboard compiles tours survey data collected  via emails sent directly to guests within 1 day post visit. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatim comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a location. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing).***"

    }

    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }

    tile button #buttonTile {
      value: "Click here to see information about guest demographics"
      navigateTo: "page_Demos"
      navigateOptions: "same_tab"

      navigateFilter: surveyDataset:filterMeasure_ToursSurvey()
    }
    label: "Voice of Guest Dashboard"
  }
  widget kpi #kpiWidget_Overall_NPS {
    label: "Overall Subsidiary NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_tours_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all tours.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Overall Subsidiary OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_tours_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Tours.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Tour(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small

    // scope reportingHierarchy {
    //   reportingHierarchy: SitesHierarchy
    //   nodes: AllData
    // }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Tour(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }


  widget headline #headlineWidget_16 {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  }
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_ToursSurvey()
      type: primary


      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_ToursSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_ToursSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_ToursSurvey()
    }
  }
  widget headline #headlineWidget_OpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_ToursSurvey()
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :PROBLEM
    }
    palette: redtogreen2ptscale

    //navigateTo: "page_Parks_Overview"
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  }
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_ToursSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small

    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_ToursSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_11 {
    label: "Recognize a Team Member?"
    hide: true
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_ToursSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget kpi #kpiWidget_Location_Value {
    label: "Tours Value"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top2percent(@reportConfig.value_qid)
      //  value: 35
      label: "Value (Top 2 Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.value_kscvc_target
    }
    infobox #infobox {
      label: "Overall Value"
      info: @reportConfig.value_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.value_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows the Value KPI for **your specific Tour(s).**  The Value KPI is based on the extent to which guests say the tour offers an ʺExtremely Goodʺ or ʺVery Goodʺ value. To see more information on Value, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.value_qid))
      label: "Average Value Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.value_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget chart #chartWidget_BookingMethod {
    label: "Booking Method"
    series #series {
      chart bar #barChart {
        showBase: true
        maxBarSize: 65
      }
      value: count(:respid)
      percentOver: "categories"
      format: noDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: noDecimalPercent
      textSize: 0
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    // chartMargin {
    //   left: 50
    // }
    layout: "horizontal"
    size: halfwidth
    category cut #cutCategory {
      value: :BOOKING_METHOD
    }
    removeEmptyCategories: true
  }
  widget comments #commentsWidget_BookingOthers {
    label: "Booking Methods - Other Specifies"

    size: small
    table: :

    sortColumn: responseColumn
    sortOrder: descending

    group question #questionGroup {
      label: "Booking Methods - Other Specify"
      filter expression #excludeBlankResponses {
        value: :BOOKING_METHOD.98$other != ""
      }
      comment: :BOOKING_METHOD.98$other
    }

    column response #responseColumn {
      sortBy: footer
      footer: :interview_start
    }

  }

  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Tours_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends"
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @NPS_Timeframe_Selector2.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector2 {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter

    }

    // scope reportingPeriod #reportingPeriodScope {
    //   period: "allData"
    // }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends"
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @OSAT_Timeframe_Selector2.selected.selectFilter
    // }

    // select #OSAT_Timeframe_Selector2 {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    // scope reportingPeriod #reportingPeriodScope {
    //   period: "allData"
    // }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "This view displays a breakdown of the performance of all locations on our key performance indicators. This provides insight on how locations perform in a relative context."


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_tours), SitesHierarchySimplified:^hierarchy) > 0

    }

    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false

    }

    column #column_current_counts {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        navigateTo: page_ToursResponses

      }

    }

    column #column_current_NPS {

      label: "NPS®"


      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        navigateTo: page_ToursResponses
       // view: comparativeStatisticView
      }
    }

    column cut #column_Promoters {
      //value: recode(@reportConfig.nps_qid, @NPScats)
      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_ToursResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends"
      // filter expression {
      //   value: @Locations_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_current_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_ToursResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }

    column #column_OSATGoal {

      label: "OSAT Goal"

      format: noDecimalNumber
      // scope reportingPeriod {
      //   period: Current
      // }
      cell {
        //value: average(numeric(SitesHierarchy:NPSTarget))
        value: parseReal(SitesHierarchySimplified:OSATTarget)
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_OSAT_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_OSAT
        other: column_OSATGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column #column_OSAT_Trends {

      // filter expression {
      //   value: @Locations_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
        }

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
      label: "Satisfaction Trends"
    }


    column #column_current_Value {
      cell #cell {
        value: top2percent(@reportConfig.value_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_ToursResponses
        navigateFilter: _isnotnull(@reportConfig.value_qid)
      }
      label: "Value (Top 2 %)"
    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget headline #headlineWidget_12 {
    label: "Key Driver Analysis By Location"
    size: large
    hide: true
    tile markdown #markdown1 {
      value: "### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

### The data below show the relationships at high levels as well as at functional levels."

//### **Please note:** These analyses require a minimum of 100 records to run; if less than 100 records are available, the report will generate an error message. If you see the message 'The accuracy of the model shown falls below the criteria specified. Please exercise caution in the use of these data.' this means that the R-squared value of the model falls below 0.5."

    }

    select #Tours_Locations_Selector {
      label: "Select a Tours Location"

      options: @valueSet_tours_locations.items

    } // end selector
  }


  widget keyDrivers #keyDriversWidget_NPS_Tours1 {
    label: "What Drives Likelihood to Recommend at " + @Tours_Locations_Selector.selectedLabel + "?"

    hide: @Tours_Locations_Selector.selected = "Tours"
    filter expression {
      value: selected(:LocationFinal, @Tours_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    //minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    minimumSampleSize: 1
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:DRILL_BOOKING.bookingsat, surveyDataset:TOURS_ELEMENTS.guidesat, surveyDataset:TOURS_ELEMENTS.sitesat

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Tours1
  widget headline #headlineWidget_9 {

    label: "Additional Key Driver Analyses for Tours locations"
    size: large
    hide: true
    select #tours_addl_keydrivers_selector {
      label: "Select an Additional Key Driver Analysis"
      options: item {
        label: "Select to see other Key Driver Analyses"
        value: 0
      },
      item {
        label: "What Drives Booking Satisfaction?"
        value: 1
      },
      item {
        label: "What Drives Tour Satisfaction?"
        value: 2
      },
      item {
        label: "What Drives Guide Satisfaction?"
        value: 3
      }


    }

    tile markdown #markdownTile_2 {
      value: "### There are several analytic views that provide us with strategic direction on what areas to promote as well as those areas that we should consider fixing . To view these, please select  an analysis from the dropdown above."
    }

  }


  widget keyDrivers #keyDriversWidget_Booking_SAT_Tours {
    label: "What Drives Booking Satisfaction at " + @Tours_Locations_Selector.selectedLabel + "?"
    hide: @tours_addl_keydrivers_selector.selected != 1

    filter expression {
      value: selected(:LocationFinal, @Tours_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:DRILL_BOOKING.bookingsat
    independentVariables: surveyDataset:DRILL_BOOKING.avail, surveyDataset:DRILL_BOOKING.info, surveyDataset:DRILL_BOOKING.communication
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_Booking_SAT_Tours
  widget keyDrivers #keyDriversWidget_Tour_SAT {
    label: "What Drives Tour Satisfaction at " + @Tours_Locations_Selector.selectedLabel + "?"
    hide: @tours_addl_keydrivers_selector.selected != 2

    filter expression {
      value: selected(:LocationFinal, @Tours_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how room features, experiences and characteristics influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT
    independentVariables: surveyDataset:TOURS_ELEMENTS.guidesat, surveyDataset:DRILL_TOURS.avail, surveyDataset:DRILL_TOURS.staff, surveyDataset:DRILL_TOURS.knowledge, surveyDataset:DRILL_TOURS.equipment
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_Tour_SAT
  widget keyDrivers #keyDriversWidget_Tour_Guide_SAT {
    label: "What Drives Guide Satisfaction at " + @Tours_Locations_Selector.selectedLabel + "?"
    hide: @tours_addl_keydrivers_selector.selected != 3

    filter expression {
      value: selected(:LocationFinal, @Tours_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation

      size: large
    }
    description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:TOURS_ELEMENTS.guidesat
    independentVariables: surveyDataset:TOURS_ELEMENTS.knowledge, surveyDataset:TOURS_ELEMENTS.toursafety, surveyDataset:TOURS_ELEMENTS.sitesat, surveyDataset:TOURS_ELEMENTS.cleanbus, surveyDataset:TOURS_ELEMENTS.lunch
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Restaurants
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  }

  widget table #tableWidget_comments {
    label: "Visitor Comments"
    size: "large"
    table: surveyDataset:

    showHeader: true
    sortOrder: descending
    sortColumn: comments

    headerNumberOfLines: 3
    stretchColumns: true
    paginationType: paging
    rowsPerPage: 100,150,250,500

    navigateTo: page_Indiv_Survey_Response
    description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response."


    select #OpenEnd_selector {
      label: "Select Question"
      options: item {
        label: "Visit Comments"
        value:  {
          selectQuestion: surveyDataset:VISIT_COMMENTS
          selectFilter: surveyDataset:VISIT_COMMENTS != ""
        }

      },
	    item {
        label: "Booking Comments"
        value:  {
          selectQuestion: surveyDataset:BOOKING_COMMENTS
          selectFilter: surveyDataset:BOOKING_COMMENTS != ""
        }

      },
	    item {
        label: "Tours Comments"
        value:  {
          selectQuestion: surveyDataset:TOURS_COMMENTS
          selectFilter: surveyDataset:TOURS_COMMENTS != ""
        }

      },
	    item {
        label: "Elements Comments"
        value:  {
          selectQuestion: surveyDataset:ELEMENTS_COMMENT
          selectFilter: surveyDataset:ELEMENTS_COMMENT != ""
        }

      },
      item {
        label: "Problem Details"
        value:  {
          selectQuestion: surveyDataset:PROBLEM_DETAIL
          selectFilter: surveyDataset:PROBLEM_DETAIL != ""
        }

      },
      item {
        label: "Team Recognition"
        value:  {
          selectQuestion: surveyDataset:RECOG_DETAIL
          selectFilter: surveyDataset:RECOG_DETAIL != ""
        }

      }      

    } // end OpenEnd_selector
    filter expression {
      value: @OpenEnd_selector.selected.selectFilter
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }


    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }


    column response #comments {
      //sortBy: comment
      header: "Location: " + surveyDataset:LocationName
      footer: @reportConfig.intvdate
     // width: 300px
      enableColumnFilter: true
      comment: @OpenEnd_selector.selected.selectQuestion

    }

    column value #LocationName {
      label: "Location"
      value: demote(SitesHierarchy:language_text, surveyDataset:)
      //value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 150px
    }


    column value #ActivityName {
      label: "Activity"
      value: :TourActivityName
      //value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 150px
    }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Rec"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    column metric #copy_of_metricColumn {
      label: "OSAT"
      value: score(@reportConfig.osat_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

    column metric #copy_of_metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

  } // end widget
  widget headline #markdownWidget_PerformanceTrends {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    }

  }

  widget dataGrid #dataGridWidget_BookingSat_Methods {
    label: "Tour Satisfaction by Booking Method"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :BOOKING_METHOD
      total: none

    }
    column #column_current_counts {

      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:BOOKING_METHOD)
        navigateTo: page_ToursResponses
       // showBase: true
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell #undefined {
        format: noDecimalPercent
        value: top1percent(:SAT)
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends"

      cell microchart {

        value: top1percent(:SAT)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_BookingSat {
    label: "Booking Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_BOOKING$field
      total: none

    }

    column #column_current_counts {
     // value: count(:SAT_EXPERIENCES$value)
      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:DRILL_BOOKING$value)
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_BOOKING$value)
        format: noDecimalPercent
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends"

      cell microchart {

        value: top1percent(:DRILL_BOOKING$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_ToursSat {
    label: "Tours Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_TOURS$field
      total: none

    }
    column #column_current_counts {

      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:DRILL_TOURS$value)
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_TOURS$value)
        format: noDecimalPercent
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends"

      cell microchart {

        value: top1percent(:DRILL_TOURS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_TourAttributesSat {
    label: "Tour Attribute Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }


    row cut {
      value: :TOURS_ELEMENTS$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:TOURS_ELEMENTS$value)
        format: noDecimalNumber
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:TOURS_ELEMENTS$value)
        format: noDecimalPercent
        navigateTo: page_ToursResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends"

      cell microchart {

        value: top1percent(:TOURS_ELEMENTS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Tours_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  modal: false
} // end page
page #page_ParksRetailFoodOverview {
  label: "Parks & Resorts - Retail / F&B"

  access rules {
    rule claim {
      name: "UserSegment"
      //value: "All", "Travel"
      value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }

  filter expression {
    value: surveyDataset:filterMeasure_DNListensParks()
    label: "DN Listens-Parks locations"
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  widget headline #headlineWidget_4 {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Parks & Resort - QR Code: Retail/F&B
### This dashboard compiles survey data collected within Parks Retail and F&B locations, collected through QR code surveys. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Trends
- Verbatims comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a single airport. 
When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }


    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_DNListensNonTravel()
    }


    label: "Voice of Guest Dashboard"
  }


  widget kpi #kpiWidget_Overall_NPS {
    label: "Parks Retail/F&B NPS®"
    size: small
    ignoreFilters: f_Location
    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all Parks Retail/F&B locations.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Parks Retail/F&B OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.osat_travel_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Parks Retail/F&B locations.**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Parks Retail/F&B location(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Parks Retail/F&B location(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Overall Satisfaction measure included in survey starting April 27, 2023"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  }
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: oneDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: primary
      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_LodgingSurvey()
    }
  }
  widget headline #headlineWidget_totalOpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small

    //     tile text #textTile0 {
    //   value: "" + @currentUser.Node
    //   fontSize: 20
    // }

    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_Recognize {
    label: "Recognize a Team Member?"
    hide: true

    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_DNListensSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"


    category cut #cutCategory {
      value: :PROBLEM

    }
    palette: redtogreen2ptscale
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  }
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Travel_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Travel_Timeframe_Selector.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Travel_Timeframe_Selector.selected.selectFilter
    // }


    // select #OSAT_Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }
    // filter expression {
    //   value: depth(SitesHierarchySimplified:^hierarchy) >= 1
    // }

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_dnlistens), SitesHierarchySimplified:^hierarchy) > 0

    }
    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row selectedFlat #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      labelStyle: nodeOnly
    //showTotal: true
    }

    column #column_current_counts {
      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
      }

    }

    column #column_current_NPS {
      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
       // target: parseReal(SitesHierarchy:NPSTarget)
        navigateTo: page_DNListensResponses
       //view: comparativeStatisticView
      }
    }

    column #column_NPSGoal {

      label: "NPS® Goal"

      format: noDecimalNumber

      cell {
        value: parseReal(SitesHierarchySimplified:NPSTarget)
        //value: average(numeric(Goals_CustomTable:nps_target))
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_NPS_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_NPS
        other: column_NPSGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column cut #column_Promoters {

      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_DNListensResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_DNListensResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }
    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

      }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs_2 {
    label: "Location KPIs (hidden)"
    size: large
    hide: true
  //ignoreFilters: reportingPeriodFilter
    removeEmptyRows: true
    description: "### For Travel Hospitality, our NPS target is 61

Note: Overall Satisfaction measure included in survey starting April 27, 2023"


    select #Locations_Timeframe_Selector {
      label: "Select Timeframe for Trends"

      options: @valueSet_date_ranges_1.items
    } // end selector
    row cut #row_2 {
      value: :LocationName
      total: "none"
    }

    column {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber

      }

    }

    column {

      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        target: @reportConfig.nps_travel_target
        navigateTo: page_DNListensResponses
        view: comparativeStatisticView
      }
    }

    column cut {

      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_DNListensResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column {
      label: "NPS® Trends"
      filter expression {
        value: @Locations_Timeframe_Selector.selected.selectFilter
      }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Locations_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

    column #column_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_DNListensResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }
    column #column_OSAT_Trends {

      filter expression {
        value: @Locations_Timeframe_Selector.selected.selectFilter
      }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Locations_Timeframe_Selector.selected.selectBreakdownBy
        }

      }

      label: "Satisfaction Trends"
    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }
  } // end widget
  // widget keyDrivers #keyDriversWidget_OSAT_Travel {
  //   label: "What Drives Guest Satisfaction?"
  //   algorithm: regression
  //   dependentVariable: @reportConfig.osat_qid
  //   independentVariables: surveyDataset:SAT_DRIVERS.quality, surveyDataset:SAT_DRIVERS.value, surveyDataset:SAT_DRIVERS.variety, surveyDataset:SAT_DRIVERS.speed, surveyDataset:SAT_DRIVERS.staff
  //   satisfactionLimit: 85
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   quadrantColors: @reportConfig.kda_quadrantColors
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_regression
  //     info: @reportConfig.kda_infobox_info_regression
  //   }
  //   description: "This analysis looks for patterns in the data to determine how guest ratings on certain experiences influence their overall satisfaction with their visit. This shows us where to target improvement initiatives."
  //   importanceLimit: 0.2
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_OSAT_Travel
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments with Text Analytics**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  }
  widget comments #commentsWidget_Dining {
    label: "Comments with Text Analytics sentiment and categories"
    size: large
    table: textAnalyticsDataset_Dining.overallScore:
    sortOrder: descending
    sortColumn: responseColumn

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000
    navigateTo: page_Indiv_Survey_Response_TA

    infobox #infobox {
      label: "Information"
      info: "This widget shows all verbatim comments, and the comment's overall sentiment or other contextual variables related to the comment. 
- Overall sentiment is measured for all the text in a comment field rather than parts of it.
- Overall sentiment ranges from -5 to 5. 0 is neutral or mixed. 
- Tags under each comment represent the topic categories associated with this comment. Tags are color-coded red for negative, yellow for neutral/mixed and green for positive. 
- Columns are filterable.
- Clicking anywhere on a comment will bring you to the Response-level results."
    }


    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: large
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: large
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
    }

    group question #questionGroup {
      label: "All Comments"
      comment: textAnalyticsDataset_Dining.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Dining.overallScore:text != ""
      }
    }
    column response #responseColumn {
      sortBy: footer
      //header: "Claim #" + surveyDataset:ClaimNbr
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta

      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "Comment Field"
      value: textAnalyticsDataset_Dining.overallScore:variable
      enableColumnFilter: true
      width: 150px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #StoreName {
      label: "Store / Restaurant"
      value: surveyDataset_TA:STORE_INFO
      enableColumnFilter: true
      //value: surveyDataset_TA:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Dining:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Dining:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 125px
    }

    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    column metric #metricColumn_NPS {
      label: "NPS"
      value: score(@reportConfig.nps_qid_ta)
      enableColumnFilter: true
      //filterable: true
      width: 125px
      align: center
      view: colorcoding
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_OSAT {
      label: "SAT"
      value: score(@reportConfig.osat_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }


    description: "**Note: To filter on Overall Sentiment, enter 3 for Positive, 2 for Neutral, 1 for Negative**
    **Note: To filter on NPS Segment, enter 3 for Promoters, 2 for Passives, 1 for Detractors**"


  } // end widget
  widget chart #TopTopics_chartWidget {

  //  label: @TANumTopics_Selector.selectedLabel + " " + @TACategoryLevels_Selector.selectedLabel + " by Volume"
    label: "Top 10 Text Analytics Topics by Volume"

    size: large
    animation: false
    gridLines: false
    legend: bottomCenter
    layout: "horizontal"
    palette: palettePosNegNueReverse

    hide: false

    filter expression {
      //value: depth(textAnalyticsDataset_Dining.model:^parent) = @TACategoryLevels_Selector.selected
      value: depth(textAnalyticsDataset_Dining.model:^parent) = 1
    }

    series #volume1 {
      label: "Mentions"
      value: textAnalyticsDataset_Dining:categoryCountTASet1()
      format: noDecimalNumber
      //navigateFilter: some(textAnalyticsDataset_Dining.categoryScore:, true, textAnalyticsDataset_Dining.categoryScore:)
      //navigateTo: dd_CategoryResultsByThemeComments
      navigateTo: dd_SentimentComments_Dining

      breakdownBy cut {
        value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      }
      percent: false
      chart bar {
        mode: stacked
        maxBarSize: 65
      }
    }
    category selectedFlat {
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
     // takeTop: @TANumTopics_Selector.selected
      takeTop: 10
      sortBy: "volume1"
      sortOrder: descending
    }


    axis secondary {
      label: "Category Sentiment"
      hide: true
    }

    axis category #categoryAxis {

      textSize: 150
      orientation: "-45"
    }
    axis primary {
      format: noDecimalNumber
    }
    navigateTo: "page_Parks_Overview"
  } // end widget
  // widget headline #headlineWidget_8 {
  //   label: "Text Analytics Sentiment Trends"
  //   size: large
  //   cardBackground: @reportConfig.selector_CardBackgroundColor


  //   select #TA_Timeframe_Selector_Dining {
  //     label: "Select a Timeframe"
  //     options: @valueSet_date_ranges.items

  //   } // end selector
  //   tile markdown #markdownTile {
  //     value: "### The section displays sentiment trends."
  //   }

  // } // end widget
  widget chart #SentimentTrends_chartWidget {
    label: "Text Analytics Sentiment Components Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
    size: large
    animation: true
    gridLines: horizontal
    legend: bottomCenter
    removeEmptyCategories: true
    hide: true
    //navigateTo: dd_SentimentComments
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Timeframe_SelectorTA1.selected.selectFilter
    // }

    infobox #infobox {
      label: "Information"
      info: "This widget shows the % distribution of overall sentiment over time. Time period break (first drop-down menu) and sentiment group base (second drop-down menu) may be selected. The distribution of the sentiment group is based on either respondents or comments for (All, positive, neutral/mixed, or negative). 
- Overall sentiment is measured for all the text in a comment field rather than parts of it. 
- Hover over the dots for more info.
- Clicking on a bar or dot will take you to the category results for that time period."
    }

    series #series_primary {
      chart bar {
        mode: "stacked100Percent"
        dataLabel: percentThenValue
        barSize: 75
        maxBarSize: 75
      }
      value: textAnalyticsDataset_Dining:overallResponseBaseTASet1()
      label: "% distribution of respondents by sentiment group"
      format: noDecimalNumber
     // format: @metric_selector.selected.cellFormat
      palette: paletteNegNeuPos
      navigateTo: dd_SentimentComments_Dining

      breakdownBy cut #cutBreakdownby {
        value: textAnalyticsDataset_Dining:responseSentimentGroup()
      }
    }

    series #series_secondary {
      value: textAnalyticsDataset_Dining:overallAverageTASet1()
      format: oneDecimalNumber
      label: "Average Sentiment"
      isSecondary: true
      chart line {
        lineWidth: 3
        dotSize: 7
        dotColorFormat: taSentimentColorDefaultFormatter
        connectNulls: true
        showDotValue: true
      }
      palette: palettePosNegNueReverse
    }


    category date #cutByDate {
      value: @reportConfig.intvdate_ta
      breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

    }

    chartMargin {
      top: 20
    }
    axis primary {
      label: "%"
      format: percentNoDecimal
      minValue: 0
      maxValue: 100
    }
    axis category {
      orientation: -45
      textSize: 75
    }
    axis secondary #secondaryAxis {
      label: "Sentiment (-5 to 5)"
      minValue: -5
      maxValue: 5
      format: noDecimalNumber
    }
    base {
      value: textAnalyticsDataset_Dining:overallResponseBaseTASet1()
      format: baseNumberFormatter
    }
    removeEmptySeries: true
  } // end widget
  widget headline #CatsAndSentiment_headlineWidget {
    label: "Text Analytics Categories & Sentiment Analysis"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #HierView_Selector {
      label: "Select a View"
      options: @valueSet_hierarchy_views.items

    } // end selector
    tile markdown #markdownTile {
      value: "###"
    }

  } // end widget
  widget dataGrid #CatsAndSentiment_HierView {
    label: "Text Analytics Categories & Sentiment - Hierarchical View"
    size: "large"

    hide: @HierView_Selector.selected != 1

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedHierarchy #comparisonRow {
      sortBy: "/percentTotalComments"
      sortOrder: descending
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:percentageOfCommentsTASet1()
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Dining:categoryCountTASet1()
        format: noDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Travel_Timeframe_Selector.selected.selectFilter
      // }
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

        }
        format: oneDecimalNumber

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Dining:categoryCount()
        extraValue: textAnalyticsDataset_Dining:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
  widget dataGrid #CatsAndSentiment_FlatView {
    label: "Text Analytics Categories & Sentiment - Flat view"
    size: "large"
    //navigateTo: dd_CategoryResultsByThemeComments

    hide: @HierView_Selector.selected != 2

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector


    row selectedFlat #comparisonRow {
      sortOrder: descending
      sortBy: "/percentTotalComments"
      reportingHierarchy: textAnalyticsDataset_Dining:categoryHierarchy_Dining
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:percentageOfCommentsTASet1()
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Dining:categoryCountTASet1()
        format: noDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Microcharts_Timeframe_Selector.selected.selectFilter
      // }
      cell microchart #cell {
        value: textAnalyticsDataset_Dining:categoryAverageTASet1()

        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy

        }
        format: oneDecimalNumber

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Dining.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Dining:categoryCount()
        extraValue: textAnalyticsDataset_Dining:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal
        //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Dining
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }

    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }
  } // end widget
  widget markdown #markdownWidget_PerformanceTrends {
    markdown: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    size: large
  }
  widget dataGrid #dataGridWidget_SatDrivers {
    label: "Satisfaction Drivers"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_DRIVERS$field
      total: none

    }
    column #column_current_counts {
      value: count(:SAT_DRIVERS$value)
      label: "Number of Responses"
      cell {
        value: count(:SAT_DRIVERS$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

    description: "Note: Variety and Value measures included in survey starting April 27, 2023.  Quality, Speed of Service, and Friendliness of Staff were included in the survey starting February 6, 2023.

Note: 'N/A' responses have been filtered out of the results below."
  } //end widget
  widget dataGrid #dataGridWidget_Sat_TimeOfDay {
    label: "Satisfaction By Time of Day"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    // sort rows {
    //   sortBy: "/Satisfaction"
    //   sortOrder: descending
    // }

    row cut {
      value: surveyDataset:TIME_OF_VISIT
      total: none

    }
    column #column_current_counts {
      value: count(surveyDataset:TIME_OF_VISIT)
      label: "Number of Responses"
      cell {
        value: count(surveyDataset:TIME_OF_VISIT)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Travel_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }


    description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023"
  } //end widget
  // widget chart #dataGridWidget_Sat_TimeOfVisit {
  //   label: "Satisfaction By Time of Visit" + " - " + @Travel_Timeframe_Selector.selectedLabel
  //   // label: @kpiselect.selected.kpiLabel + " Trends"   
  //   palette: multicolors1_palette
  //  // ignoreFilters: reportingPeriodFilter

  //   // select #TimeofDay_Timeframe_Selector {
  //   //   label: "Select Timeframe"

  //   //   options: @valueSet_date_ranges_1.items

  //   // } // end selector
  //   size: halfwidth

  //   legend: bottomCenter
  //   chartMargin {
  //     top: 20
  //     bottom: 75
  //     right: 25
  //   }

  //   series #series {
  //     chart line {
  //       showDotValue: false

  //     }

  //     value: top1percent(@reportConfig.osat_qid)
  //     format: oneDecimalPercent

  //     isSecondary: false
  //     breakdownBy cut {
  //       value: surveyDataset:TIME_OF_VISIT

  //     }
  //   }

  //   category date #dateCategory {
  //     value: @reportConfig.intvdate
  //     breakdownBy: @Travel_Timeframe_Selector.selected.selectBreakdownBy
  //     label: "Interview date"
  //     //format: dateDefaultFormatter
  //   }


  //   axis category #categoryAxis {
  //     orientation: "-45"
  //     format: noDecimalPercent

  //   }
  //   axis primary #primaryAxis {
  //        //  format: metricsItemMetricDefaultFormatter
  //     format: noDecimalPercent
  //     label: "% Very Satisfied"
  //     minValue: 50
  //     maxValue: 100
  //   }
  //   axis secondary #secondaryAxis {
  //     hide: true
  //     label: "% Response"
  //     format: noDecimalPercent
  //     minValue: 0
  //     maxValue: 100
  //   }


  //   base #base {
  //     value: count(@reportConfig.osat_qid)
  //     format: baseNumberFormatter
  //   }
  //   removeEmptyCategories: true
  //   removeEmptySeries: true
  // } // end widget
} // end page
page #page_Gaming_Overview {
  label: "Gaming"
  //hide: true
  modal: false

  access rules {
    rule claim {
      name: "UserSegment"
      value: "All", "Gaming"
      //value: "Test"
    }
  }


  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_GamingSurvey()
    label: "Gaming survey Only"
  }


  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }


  layoutArea toolbar {
    filter multiselect #f_LoyaltyTier {
      label: "Loyalty Tier"
      optionsFrom: :rank_description
    }
  }
  widget headline #headlineWidget_Gaming_Overview {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Gaming  Dashboard
### This dashboard compiles gaming survey data collected  via emails sent directly to guests within 1 day post visit. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatim comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a location. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }

    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }

    tile button #buttonTile {
      value: "Click here to see information about guest demographics"
      navigateTo: "page_Demos_Gaming"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_GamingSurvey()
    }
    label: "Voice of Guest Dashboard"
  }
  widget kpi #kpiWidget_Overall_NPS {
    label: "Overall Subsidiary NPS®"
    size: small
    ignoreFilters: f_Location

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_ExcludeAustraliaLocations()
      label: "Exclude Australia locations"
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.nps_gaming_target
    }
    infobox #infobox {
      label: "NPS®"
      info: "The Net Promoter Score®, or NPS®, is a way of assessing the level of loyalty that a customer has toward an organization. We first ask a question about the customer's likelihood to recommend us:

ʺBased on your recent visit, on a scale from 0 to 10, how likely are you to recommend this location to a friend or family member? ʺ

Customers rating a 9 or 10 are called Promoters - these are the most favorable customers; on the other end of the spectrum, we have Detractors - those who rate from 0 to 6 on the scale. Customers rating 7 or 8 are put into a category called Passives.

To calculate the NPS®, we take the percentage of Promoters and subtract the percentage of Detractors. This means that NPS can fall on a scale between -100 (no Promoters) to 100 (all Promoters).

What should we do with this information? It can help with our efforts to act on customer insight - for example, Promoters are customers who are more likely to buy more (or different) products; they can also be great references. Detractors, on the other hand, often provide insight on areas of friction that we should consider Fixing."
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **all Gaming locations.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above.

Note: Australia locations have been excluded on this widget."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }

  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Overall Subsidiary OSAT"
    size: small
    ignoreFilters: f_Location

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_ExcludeAustraliaLocations()
      label: "Exclude Australia locations"
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_gaming_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **all Gaming locations.**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.

Note: Australia locations have been excluded on this widget.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Gaming location(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small

    // scope reportingHierarchy {
    //   reportingHierarchy: SitesHierarchy
    //   nodes: AllData
    // }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Gaming location(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  } // end widget
  widget markdown #headlineWidget_NPS_Cats {
    pageBreak: true
    size: large
    markdown: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
  }
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_GamingSurvey()
      type: primary


      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_GamingSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_GamingSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_GamingSurvey()
    }
  }
  widget headline #headlineWidget_OpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_GamingSurvey()
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :PROBLEM
    }
    palette: redtogreen2ptscale

    navigateTo: "page_Parks_Overview"
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  } // end widget
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_GamingSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  } // end widget
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small


    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_GamingSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_Recognize {
    label: "Recognize a Team Member?"
    hide: true
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_GamingSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Gaming_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @NPS_Timeframe_Selector_Gaming.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector_Gaming {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }


      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter

    }

    // scope reportingPeriod #reportingPeriodScope {
    //   period: "allData"
    // }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @OSAT_Timeframe_Selector_Gaming.selected.selectFilter
    // }

    // select #OSAT_Timeframe_Selector_Gaming {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    // scope reportingPeriod #reportingPeriodScope {
    //   period: "allData"
    // }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "### This view displays a breakdown of the performance of all locations on our key performance indicators. This provides insight on how locations perform in a relative context.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"


    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }


    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_gaming), SitesHierarchySimplified:^hierarchy) > 0

    }

    // select #Locations_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_current_counts {
      label: "n"
      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }

    }

    column #column_current_NPS {

      label: "NPS®"

      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        navigateTo: page_GamingResponses
       // view: comparativeStatisticView
      }
    }

    column #column_NPSGoal {

      label: "NPS® Goal"

      format: noDecimalNumber
      // scope reportingPeriod {
      //   period: Current
      // }
      cell {
        //for any locaitons without a target, set target to "TBD" in the table
        value: parseReal(SitesHierarchySimplified:NPSTarget)

        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_NPS_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_NPS
        other: column_NPSGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column cut #column_Promoters {
      //value: recode(@reportConfig.nps_qid, @NPScats)
      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        navigateTo: page_GamingResponses
        navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }


    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column {
      label: "NPS® Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Locations_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_current_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        navigateTo: page_GamingResponses
        navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }

    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Locations_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        }

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget headline #headlineWidget_KDAs_Location {
    label: "Key Driver Analysis By Location"
    size: large

    tile markdown #markdown1 {
      value: "### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

### The data below show the relationships at high levels as well as at functional levels. "

    }

    select #Gaming_Locations_Selector {
      label: "Select a Gaming Location"

      options: @valueSet_gaming_locations.items

    } // end selector
  }
  widget keyDrivers #keyDriversWidget_NPS_Gaming1 {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among casino visitors?"

  //attributes removed for this KDA: lodging
  //this kda applies to following locations:
    //SL	Southland Casino
    //WI	Wheeling Island - Casino - Racetrack

    hide: @Gaming_Locations_Selector.selected.selectCode != "SL" AND @Gaming_Locations_Selector.selected.selectCode != "WI"

    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.buffet, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.pokerroom, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots, surveyDataset:SAT_GAMING.tablegames


    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming1
  widget keyDrivers #keyDriversWidget_NPS_Gaming2 {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among casino visitors?"

  //attributes removed for this KDA: lodging, buffet
  //this kda applies to following locations:
    //BB	Gate City Casino (formerly Boston Billiards)
    //DB	Daytona Beach Racing and Card Club
    //OC	Orange City Racing and Card Club
    //MB	Mindil Beach Casino Resort
    //MG	Mardi Gras Casino & Resort

    hide: @Gaming_Locations_Selector.selected.selectCode != "BB" AND @Gaming_Locations_Selector.selected.selectCode != "DB" AND @Gaming_Locations_Selector.selected.selectCode != "OC" AND @Gaming_Locations_Selector.selected.selectCode != "MBCR" AND @Gaming_Locations_Selector.selected.selectCode != "MG"
    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    // minimumSampleSize: 1  
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.pokerroom, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots, surveyDataset:SAT_GAMING.tablegames

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming2
  widget keyDrivers #keyDriversWidget_NPS_Gaming3 {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among casino visitors?"

  //attributes removed for this KDA: lodging, buffet, poker room, tablegames
  //this kda applies to following locations:
    //HB	Hamburg Gaming

    hide: @Gaming_Locations_Selector.selected.selectCode != "HB"

    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming3
  widget keyDrivers #keyDriversWidget_NPS_Gaming4 {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among casino visitors?"

  //attributes removed for this KDA: lodging, buffet, poker room, tablegames
  //this kda applies to following locations:
    //MVG	Miami Valley Gaming & Racing

    hide: @Gaming_Locations_Selector.selected.selectCode != "MVG"

    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming4
  widget keyDrivers #keyDriversWidget_NPS_Gaming5 {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among casino visitors?"

  //attributes removed for this KDA: lodging, poker room, tablegames
  //this kda applies to following locations:
    //FL	Finger Lakes Gaming & Racetrack

    hide: @Gaming_Locations_Selector.selected.selectCode != "FL"

    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    // minimumSampleSize: 1  
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.buffet, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming5
  widget keyDrivers #keyDriversWidget_NPS_Gaming7 {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among casino visitors?"

  //attributes removed for this KDA: lodging, bars, buffet, pokerroom, tablegames
  //this kda applies to following locations:
    //TK	Catawba Two Kings Casino

    hide: @Gaming_Locations_Selector.selected.selectCode != "TK"

    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.buffet, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming7
  widget keyDrivers #keyDriversWidget_NPS_Gaming_MG_hotel {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among hotel guests?"

  //attributes removed for this KDA: buffet
  //this kda applies to following locations:
    //7689	Mardi Gras Casino & Resort Hotel

    hide: @Gaming_Locations_Selector.selected.selectCode != "MG"

    filter expression {
      //7689	Mardi Gras Casino & Resort Hotel
      value: selected(:LocationFinal, "7689")

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "" + @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.lodging, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.pokerroom, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots, surveyDataset:SAT_GAMING.tablegames

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming_MG_hotel
  widget keyDrivers #keyDriversWidget_NPS_Gaming_SL_hotel {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among hotel guests?"

  //attributes removed for this KDA: none
  //this kda applies to following locations:
    //38344	Southland Casino Hotel

    hide: @Gaming_Locations_Selector.selected.selectCode != "SL"

    filter expression {
      //7689	Mardi Gras Casino & Resort Hotel
      value: selected(:LocationFinal, "38344")

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.buffet, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.lodging, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.pokerroom, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots, surveyDataset:SAT_GAMING.tablegames

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming_SL_hotel
  widget keyDrivers #keyDriversWidget_NPS_Gaming_WI_hotel {
    label: "What Drives Likelihood to Recommend at " + @Gaming_Locations_Selector.selectedLabel + " among hotel guests?"

  //attributes removed for this KDA: bars
  //this kda applies to following locations:
    //51559	Wheeling Island Hotel - Casino - Racetrack

    hide: @Gaming_Locations_Selector.selected.selectCode != "WI"

    filter expression {
      //51559	Wheeling Island Hotel - Casino - Racetrack
      value: selected(:LocationFinal, "51559")

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    //algorithm: regression
    algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      // label: @reportConfig.kda_infobox_label_regression
      // info: @reportConfig.kda_infobox_info_regression

      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.buffet, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.lodging, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.pokerroom, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.slots, surveyDataset:SAT_GAMING.tablegames

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Gaming_SL_hotel
  widget headline #headlineWidget_KDAs_Location_Addtl {

    label: "Additional Key Driver Analyses for " + @Gaming_Locations_Selector.selectedLabel + ""
    size: large

    select #gaming_addl_keydrivers_selector {
      label: "Select an Additional Key Driver Analysis"
      options: item {
        label: "Select to see other Key Driver Analyses"
        value: 0
      },
      item {
        label: "What Drives Satisfaction with Gaming?"
        value: 1
      },
      item {
        label: "What Drives Satisfaction with Slots/Gaming Machines?"
        value: 2
      },
      item {
        label: "What Drives Satisfaction with Table Games?"
        value: 3
      },
      item {
        label: "What Drives Satisfaction with Lodging?"
        value: 4
      },
      item {
        label: "How Do Room Features Impact Lodging Satisfaction?"
        value: 5
      },
      item {
        label: "What Drives Restaurant Satisfaction?"
        value: 6
      },
      item {
        label: "What Drives Buffet Satisfaction?"
        value: 7
      },
      item {
        label: "What Drives Bar Satisfaction?"
        value: 8
      }
    }

    tile markdown #markdownTile_2 {
      value: "### There are several analytic views that provide us with strategic direction on what areas to promote as well as those areas that we should consider fixing . To view these, please select  an analysis from the dropdown above."
    }

  }
  widget keyDrivers #keyDriversWidget_SAT_Gaming {
    label: "What Drives Satisfaction with Gaming at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 1
    filter expression {
      value: @Gaming_Locations_Selector.selected.selectFilter

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT
    independentVariables: surveyDataset:SAT_DRIVERS.cleanliness, surveyDataset:SAT_DRIVERS.knowledge, surveyDataset:SAT_DRIVERS.speed, surveyDataset:SAT_DRIVERS.safety, surveyDataset:SAT_DRIVERS.staff, surveyDataset:SAT_DRIVERS.valet
    warningText: @reportConfig.kda_warningText
 //   rSquaredLimit: 0.5
  } // end widget keyDriversWidget_SAT_Gaming
  widget keyDrivers #keyDriversWidget_SAT_Slots {
    label: "What Drives Satisfaction with Slots/Gaming Machines at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 2
    filter expression {
      value: @Gaming_Locations_Selector.selected.selectFilter

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall gaming satisfaction. This shows us where to target improvement in our gaming processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_GAMING.slots
    independentVariables: surveyDataset:DRILL_SLOTS.avail, surveyDataset:DRILL_SLOTS.selection
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Slots
  widget keyDrivers #keyDriversWidget_SAT_TableGames {
    label: "What Drives Satisfaction with Table Games at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 3
    filter expression {
      value: @Gaming_Locations_Selector.selected.selectFilter

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall gaming satisfaction. This shows us where to target improvement in our gaming processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_GAMING.tablegames
    independentVariables: surveyDataset:DRILL_TABLEGAMES.avail, surveyDataset:DRILL_TABLEGAMES.betting, surveyDataset:DRILL_TABLEGAMES.selection, surveyDataset:DRILL_TABLEGAMES.staff
    warningText: @reportConfig.kda_warningText
    //rSquaredLimit: 0.9
  } // end widget keyDriversWidget_SAT_TableGames
  widget keyDrivers #keyDriversWidget_SAT_Lodging {
    label: "What Drives Satisfaction with Lodging at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 4
    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectHotelCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall gaming satisfaction. This shows us where to target improvement in our gaming processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT_GAMING.lodging
    independentVariables: surveyDataset:DRILL_LODGING.ease, surveyDataset:DRILL_LODGING.accuracy, surveyDataset:DRILL_LODGING.arrival, surveyDataset:DRILL_LODGING.cleanliness, surveyDataset:DRILL_LODGING.avail, surveyDataset:DRILL_LODGING.departure, surveyDataset:DRILL_LODGING.service
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Lodging
  widget keyDrivers #keyDriversWidget_SAT_Room {
    label: "How Do Room Features Impact Lodging Satisfaction at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 5
    filter expression {
      value: selected(:LocationFinal, @Gaming_Locations_Selector.selected.selectHotelCode)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how room features, experiences and characteristics influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT_GAMING.lodging
    independentVariables: surveyDataset:DRILL_ROOM.ac, surveyDataset:DRILL_ROOM.bathclean, surveyDataset:DRILL_ROOM.bathfeatures, surveyDataset:DRILL_ROOM.bed, surveyDataset:DRILL_ROOM.cleanliness, surveyDataset:DRILL_ROOM.quiet, surveyDataset:DRILL_ROOM.wifi, surveyDataset:DRILL_ROOM.bathamenities, surveyDataset:DRILL_ROOM.smell, surveyDataset:DRILL_ROOM.furnishings
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Room
  widget keyDrivers #keyDriversWidget_SAT_Restaurants {
    label: "What Drives Restaurant Satisfaction at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 6
    filter expression {
      value: @Gaming_Locations_Selector.selected.selectFilter

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    select #catfilter {
      label: "Filter by Meal Rated"
      mode: multi

      options: @categorySet_meal_rated.items
    }
    filter expression {
      value: selected(:MEAL_RATED, @catfilter.selected)
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation

      size: large
    }
    description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_GAMING.restaurants
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.quality, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.variety
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Restaurants
  widget keyDrivers #keyDriversWidget_SAT_Buffet {
    label: "What Drives Buffet Satisfaction at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 7
    filter expression {
      value: @Gaming_Locations_Selector.selected.selectFilter

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the buffet influence their overall buffet satisfaction. This shows us where to target improvement in our buffet processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_GAMING.buffet
    independentVariables: surveyDataset:DRILL_BUFFET.cleanliness, surveyDataset:DRILL_BUFFET.quality, surveyDataset:DRILL_BUFFET.stock, surveyDataset:DRILL_BUFFET.taste, surveyDataset:DRILL_BUFFET.temperature, surveyDataset:DRILL_BUFFET.value, surveyDataset:DRILL_BUFFET.variety
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Buffet
  widget keyDrivers #keyDriversWidget_SAT_Bars {
    label: "What Drives Bar Satisfaction at " + @Gaming_Locations_Selector.selectedLabel + "?"
    hide: @gaming_addl_keydrivers_selector.selected != 8
    filter expression {
      value: @Gaming_Locations_Selector.selected.selectFilter

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 86
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the bar influence their overall bar satisfaction. This shows us where to target improvement in our bar processes and experiences."
    importanceLimit: 0.25
    dependentVariable: surveyDataset:SAT_GAMING.bars
    independentVariables: surveyDataset:DRILL_GAME_DRINK.speed, surveyDataset:DRILL_GAME_DRINK.taste, surveyDataset:DRILL_GAME_DRINK.value
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Bars
  widget headline #headlineWidget_14 {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments with Text Analytics**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  }
  widget comments #commentsWidget {
    label: "Comments with Text Analytics sentiment and categories"
    size: large
    table: textAnalyticsDataset_Gaming.overallScore:
    sortOrder: descending
    sortColumn: responseColumn

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response_TA

    infobox #infobox {
      label: "Information"
      info: "This widget shows all verbatim comments, and the comment's overall sentiment or other contextual variables related to the comment. 
- Overall sentiment is measured for all the text in a comment field rather than parts of it.
- Overall sentiment ranges from -5 to 5. 0 is neutral or mixed. 
- Tags under each comment represent the topic categories associated with this comment. Tags are color-coded red for negative, yellow for neutral/mixed and green for positive. 
- Columns are filterable.
- Clicking anywhere on a comment will bring you to the Response-level results."
    }


    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
      fontSize: medium
    }

    group question #questionGroup {
      label: "All Comments"
      comment: textAnalyticsDataset_Gaming.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Gaming.overallScore:text != ""
      }
    }
    column response #responseColumn {
      sortBy: footer
      //header: "Claim #" + surveyDataset:ClaimNbr
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta

      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "Comment Field"
      value: textAnalyticsDataset_Gaming.overallScore:variable
      enableColumnFilter: true
      width: 150px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #LoyaltyTier {
      label: "Loyalty Tier"
      value: surveyDataset:rank_description
      //value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 100px
    }

    column metric #metricColumn {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Gaming:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Lodging:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 125px
    }

    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    column metric #metricColumn_NPS {
      label: "NPS"
      value: score(@reportConfig.nps_qid_ta)
      enableColumnFilter: true
      //filterable: true
      width: 125px
      align: center
      view: colorcoding
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_OSAT {
      label: "SAT"
      value: score(@reportConfig.osat_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }

    column metric #metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false //hides from screen but is exported
    }



    description: "**Note: To filter on Overall Sentiment, enter 3 for Positive, 2 for Neutral, 1 for Negative**
    **Note: To filter on NPS Segment, enter 3 for Promoters, 2 for Passives, 1 for Detractors**"


  } // end widget
  widget chart #TopTopics_chartWidget {

  //  label: @TANumTopics_Selector.selectedLabel + " " + @TACategoryLevels_Selector.selectedLabel + " by Volume"
    label: "Top 10 Text Analytics Topics by Volume"

    size: large
    animation: false
    gridLines: false
    legend: bottomCenter
    layout: "horizontal"
    palette: palettePosNegNueReverse

    hide: false

    filter expression {
      //value: depth(textAnalyticsDataset_Lodging.model:^parent) = @TACategoryLevels_Selector.selected
      value: depth(textAnalyticsDataset_Gaming.model:^parent) = 2
    }

    series #volume1 {
      label: "Mentions"
      value: textAnalyticsDataset_Gaming:categoryCountTASet1()
      format: noDecimalNumber
      //navigateFilter: some(textAnalyticsDataset_Lodging.categoryScore:, true, textAnalyticsDataset_Lodging.categoryScore:)
      //navigateTo: dd_CategoryResultsByThemeComments
      navigateTo: dd_SentimentComments_Gaming

      breakdownBy cut {
        value: textAnalyticsDataset_Gaming.categoryScore:categorySentimentGroup
      }
      percent: false
      chart bar {
        mode: stacked
        maxBarSize: 65
      }
    }
    category selectedFlat {
      reportingHierarchy: textAnalyticsDataset_Gaming:categoryHierarchy_Gaming
     // takeTop: @TANumTopics_Selector.selected
      takeTop: 10
      sortBy: "volume1"
      sortOrder: descending
    }


    axis secondary {
      label: "Category Sentiment"
      hide: true
    }

    axis category #categoryAxis {

      textSize: 100
      orientation: "-45"
    }
    axis primary {
      format: noDecimalNumber
    }
    navigateTo: "page_Gaming_Overview"
  } // end widget
  widget chart #SentimentTrends_chartWidget {
    label: "Text Analytics Sentiment Components Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel
    size: large
    animation: true
    gridLines: horizontal
    legend: bottomCenter
    removeEmptyCategories: true
    //navigateTo: dd_SentimentComments
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @Timeframe_SelectorTA1.selected.selectFilter
    // }

    infobox #infobox {
      label: "Information"
      info: "This widget shows the % distribution of overall sentiment over time. Time period break (first drop-down menu) and sentiment group base (second drop-down menu) may be selected. The distribution of the sentiment group is based on either respondents or comments for (All, positive, neutral/mixed, or negative). 
- Overall sentiment is measured for all the text in a comment field rather than parts of it. 
- Hover over the dots for more info.
- Clicking on a bar or dot will take you to the category results for that time period."
    }

    series #series_primary {
      chart bar {
        mode: "stacked100Percent"
        dataLabel: percentThenValue
        barSize: 75
        maxBarSize: 75
      }
      value: textAnalyticsDataset_Gaming:overallResponseBaseTASet1()
      label: "% distribution of respondents by sentiment group"
      format: noDecimalNumber
     // format: @metric_selector.selected.cellFormat
      palette: paletteNegNeuPos
      navigateTo: dd_SentimentComments_Gaming

      breakdownBy cut #cutBreakdownby {
        value: textAnalyticsDataset_Gaming:responseSentimentGroup()
      }
    }

    series #series_secondary {
      value: textAnalyticsDataset_Gaming:overallAverageTASet1()
      format: oneDecimalNumber
      label: "Average Sentiment"
      isSecondary: true
      chart line {
        lineWidth: 3
        dotSize: 7
        dotColorFormat: taSentimentColorDefaultFormatter
        connectNulls: true
        showDotValue: true
      }
      palette: palettePosNegNueReverse
    }


    category date #cutByDate {
      value: @reportConfig.intvdate_ta
      breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    chartMargin {
      top: 20
    }
    axis primary {
      label: "%"
      format: percentNoDecimal
      minValue: 0
      maxValue: 100
    }
    axis category {
      orientation: -45
      textSize: 75
    }
    axis secondary #secondaryAxis {
      label: "Sentiment (-5 to 5)"
      minValue: -5
      maxValue: 5
      format: noDecimalNumber
    }
    base {
      value: textAnalyticsDataset_Gaming:overallResponseBaseTASet1()
      format: baseNumberFormatter
    }
    removeEmptySeries: true
  } // end widget
  widget headline #CatsAndSentiment_headlineWidget {
    label: "Text Analytics Categories & Sentiment Analysis"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #HierView_Selector {
      label: "Select a View"
      options: @valueSet_hierarchy_views.items

    } // end selector
    tile markdown #markdownTile {
      value: "###"
    }

  } // end widget
  widget dataGrid #CatsAndSentiment_HierView {
    label: "Text Analytics Categories & Sentiment - Hierarchical View"
    size: "large"

    hide: @HierView_Selector.selected != 1

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedHierarchy #comparisonRow {
      sortBy: "/percentTotalComments"
      sortOrder: descending
      reportingHierarchy: textAnalyticsDataset_Gaming:categoryHierarchy_Gaming
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Gaming:percentageOfCommentsTASet1()
        format: percentNoDecimal
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Gaming
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Gaming:categoryCountTASet1()
        format: noDecimalNumber

        navigateTo: dd_SentimentComments_Gaming
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Gaming:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber

        navigateTo: dd_SentimentComments_Gaming
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel
      filter expression {
        value: @Gaming_Timeframe_Selector.selected.selectFilter
      }
      cell microchart #cell {
        value: textAnalyticsDataset_Gaming:categoryAverageTASet1()
        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
          align: true
          //start: "-4 quarter"

        }
        format: oneDecimalNumber

      }

    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Gaming.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Gaming:categoryCount()
        extraValue: textAnalyticsDataset_Gaming:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal

        navigateTo: dd_SentimentComments_Gaming
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
  widget dataGrid #CatsAndSentiment_FlatView {
    label: "Text Analytics Categories & Sentiment - Flat view"
    size: "large"


    hide: @HierView_Selector.selected != 2

    // select #Microcharts_Timeframe_Selector {
    //   label: "Select Timeframe for Trends"

    //   options: @valueSet_date_ranges.items
    // } // end selector
    infobox #infobox {
      label: "Information"
      info: " This widget shows a detailed table view of the nested category taxonomy, category volume, and category sentiment. Category sentiment is measured for the section of the comment field which aligns to the model's category definitions.  
- Each row shows the results of each category , with the ability  to drill down to see results of sub-categories, where a sub-category is available.
- In the first column you have the ability to drill down and see sub categories within a model name.  
- Clicking on individual cells go to the comments for that cell.
- Please select a specific category or categories in the filter on the left to limit the view."
    }

    row selectedFlat #comparisonRow {
      sortOrder: descending
      sortBy: "/percentTotalComments"
      reportingHierarchy: textAnalyticsDataset_Gaming:categoryHierarchy_Gaming
      showTotal: false
    }
    column #percentTotalComments {
      label: "% of Total Comments"
      cell microchart #cell {
        value: textAnalyticsDataset_Gaming:percentageOfCommentsTASet1()
        format: percentNoDecimal
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Gaming
        microchart bar #barMicrochart {
          colorFormat: dropOffDefaultFormatter
          valuePosition: outer
          min: 0
          max: 100
        }
      }
    }
    column #numberComments {
      label: "# Comments"
      cell #cell {
        value: textAnalyticsDataset_Gaming:categoryCountTASet1()
        format: noDecimalNumber
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Gaming
      }
    }
    column #avgSentiment {
      label: "Avg. Sentiment"

      cell #cell {
        value: textAnalyticsDataset_Gaming:categoryAverageTASet1()
        view: sentimentView
        format: oneDecimalNumber
      //navigateTo: dd_CategoryResultsByThemeComments
        navigateTo: dd_SentimentComments_Gaming
      }
    }
    column #sentimentTrend {
      label: "Sentiment Trends"

      cell microchart #cell {
        value: textAnalyticsDataset_Gaming:categoryAverageTASet1()

        useOnlyExistingColumns: true

        microchart line #barMicrochart {
          min: auto
          max: auto
          color: #004d63
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate_ta
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
          align: true
          //start: "-4 quarter"
        }
        format: oneDecimalNumber

      }

    }
    column cut #percentCommentsCategory {
      label: "% of Comments Within Category"
      value: textAnalyticsDataset_Gaming.categoryScore:categorySentimentGroup
      total: "none"
      showLabel: true
      cell columnPercentage #cell {
        value: textAnalyticsDataset_Gaming:categoryCount()
        extraValue: textAnalyticsDataset_Gaming:categoryCount()
        extraValueFormat: noDecimalNumber
        format: percentNoDecimal

        navigateTo: dd_SentimentComments_Gaming
      }
    }
    view comparativeStatistic #sentimentView {
      backgroundColorFormatter: taSentimentColorDefaultFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }
  } // end widget
//   widget markdown #headlineWidget_Comments {
//     markdown: "## **Guest Comments**

// ### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

// ### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
//     size: large
//   }
//   widget table #tableWidget_Comments {
//     label: "Visitor Comments"
//     size: "large"
//     table: surveyDataset:

//     showHeader: true
//     sortOrder: descending
//     sortColumn: comments

//     headerNumberOfLines: 3
//     stretchColumns: true

//     paginationType: paging
//     rowsPerPage: 100, 250, 500, 1000


//     navigateTo: page_Indiv_Survey_Response
//     description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response."


//     select #OpenEnd_selector {
//       label: "Select Question"
//       options: item {
//         label: "Visit Comments"
//         value:  {
//           selectQuestion: surveyDataset:VISIT_COMMENTS
//           selectFilter: surveyDataset:VISIT_COMMENTS != ""
//         }

//       },
// 	    item {
//         label: "Lodging Comments"
//         value:  {
//           selectQuestion: surveyDataset:LODGING_COMMENTS
//           selectFilter: surveyDataset:LODGING_COMMENTS != ""
//         }

//       },
// 	    item {
//         label: "Restaurant/Buffet Comments"
//         value:  {
//           selectQuestion: surveyDataset:RESTAURANT_COMMENTS
//           selectFilter: surveyDataset:RESTAURANT_COMMENTS != ""
//         }

//       },
//       item {
//         label: "Problem Details"
//         value:  {
//           selectQuestion: surveyDataset:PROBLEM_DETAIL
//           selectFilter: surveyDataset:PROBLEM_DETAIL != ""
//         }

//       },
//       item {
//         label: "Team Recognition"
//         value:  {
//           selectQuestion: surveyDataset:RECOG_DETAIL
//           selectFilter: surveyDataset:RECOG_DETAIL != ""
//         }

//       }    

//     } // end OpenEnd_selector
//     filter expression {
//       value: @OpenEnd_selector.selected.selectFilter
//     }

//     view metric #viewnpssegment {
//       backgroundColorFormatter: sentimentindicator2a //backgroundColor 
//       valueColorFormatter: sentimentindicator2text //textColors
//       fontSize: medium
//     }


//     view metric #colorcoding_11pt {
//       backgroundColorFormatter: sentimentindicator1 //backgroundColor 
//       valueColorFormatter: sentimentindicator1text //textColors
//       fontSize: medium
//     }

//     view metric #colorcoding_5pt {
//       backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
//       valueColorFormatter: sentimentindicator_text_5pt //textColors
//       fontSize: medium
//     }


//     column response #comments {
//       //sortBy: comment
//       header: "Location: " + surveyDataset:LocationName
//       footer: @reportConfig.intvdate
//      // width: 300px
//       enableColumnFilter: true
//       comment: @OpenEnd_selector.selected.selectQuestion

//     }


//     // column value #SurveyName {
//     //   label: "Survey"
//     //   value: surveyDataset:survey_name
//     //   enableColumnFilter: true
//     //   align: center
//     //   width: 150px

//     // }


//     column value #LocationName {
//       label: "Location"
//       value: demote(SitesHierarchy:language_text, surveyDataset:)
//       //value: surveyDataset:LocationName
//       enableColumnFilter: true
//       //value: surveyDataset:SitesHierarchy
//       width: 200px
//     }

//     column value #LoyaltyTier {
//       label: "Loyalty Tier"
//       value: surveyDataset:rank_description
//       //value: surveyDataset:LocationName
//       enableColumnFilter: true
//       //value: surveyDataset:SitesHierarchy
//       width: 100px
//     }

//     column metric #metricColumn_1 {
//       label: "NPS Segment"
//       value: score(surveyDataset:NPSVal)
//       format: npssegmentindicatortextValue2
//       target: 9
//       view: viewnpssegment
//       width: 100px
//       align: center
//       enableColumnFilter: true
//     }

//     column metric #metricColumn {
//       label: "Likely to Rec"
//       value: @reportConfig.nps_qid
//       enableColumnFilter: true
//       width: 100px
//       align: center
//       view: colorcoding_11pt

//     }
//     column metric #copy_of_metricColumn {
//       label: "OSAT"
//       value: score(@reportConfig.osat_qid)
//       enableColumnFilter: true
//       width: 100px
//       align: center
//       view: colorcoding_5pt

//     }

//   } // end widget
  widget markdown #markdownWidget_PerformanceTrends {
    markdown: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of gaming. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    size: large
  }
  widget dataGrid #dataGridWidget_SatDrivers {
    label: "Satisfaction Drivers"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_DRIVERS$field
      total: none

    }
    column #column_current_counts {
      value: count(:SAT_DRIVERS$value)
      label: "Number of Responses"
      cell {
        value: count(:SAT_DRIVERS$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_GamingSat {
    label: "Gaming Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_GAMING$field
      total: none

    }
    column #column_current_counts {
      value: count(:SAT_GAMING$value)
      label: "Number of Responses"
      cell {
        value: count(:SAT_GAMING$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:SAT_GAMING$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_GAMING$value)
        format: noDecimalPercent

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_SlotsSat {
    label: "Slots Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_SLOTS$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_SLOTS$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_SLOTS$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_SLOTS$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_SLOTS$value)
        format: noDecimalPercent

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_TableGamesSat {
    label: "Table Games Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_TABLEGAMES$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_TABLEGAMES$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_TABLEGAMES$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_TABLEGAMES$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_TABLEGAMES$value)
        format: noDecimalPercent

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_DrinkSat {
    label: "Drink Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_GAME_DRINK$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_GAME_DRINK$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_GAME_DRINK$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_GAME_DRINK$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_GAME_DRINK$value)
        format: noDecimalPercent

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_LodgingSat {
    label: "Lodging Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_LODGING$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_LODGING$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_LODGING$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        extraValue: count(:DRILL_LODGING$value)
        extraValueFormat: noDecimalNumber
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_RoomSat {
    label: "Room Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_ROOM$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_ROOM$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_ROOM$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_BuffetSat {
    label: "Buffet Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_BUFFET$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_BUFFET$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_BUFFET$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_BUFFET$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_RestaurantSat {
    label: "Restaurant Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    select #catfilter {
      label: "Filter by Meal Rated"
      mode: multi

      options: @categorySet_meal_rated.items
    }
    filter expression {
      value: selected(:MEAL_RATED, @catfilter.selected)
    }

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_RESTAURANT$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_RESTAURANT$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_RESTAURANT$value)
        format: noDecimalNumber
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        navigateTo: page_GamingResponses
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_Sat_LoyaltyTier {
    label: "Satisfaction By Loyalty Tier"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    // sort rows {
    //   sortBy: "/Satisfaction"
    //   sortOrder: descending
    // }

    row cut {
      value: surveyDataset:LoyaltyTiers
      total: none
    }


    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent
        extraValue: count(@reportConfig.osat_qid)
        extraValueFormat: noDecimalNumber
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

    column #column_Responses_Trends {
      label: "Number of Responses Trends" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: count(@reportConfig.osat_qid)
        format: noDecimalNumber
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

    //description: "Note: Overall Satisfaction measure included in survey starting April 27, 2023"
  } //end widget
  widget dataGrid #dataGridWidget_SatByLoyaltyTier {
    label: "Satisfaction By Loyalty Tier"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    removeEmptyColumns: true
    description: ""

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }

    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row cut {
      value: surveyDataset:LocationName
      showTotal: false
    }


    column #column_OSAT {
      label: "% Satisfied (Top Box)"
      column cut {
        total: none
        value: surveyDataset:LoyaltyTiers

        cell #cell {
          value: top1percent(@reportConfig.osat_qid)
          format: noDecimalPercent
          extraValue: count(@reportConfig.osat_qid)
          extraValueFormat: noDecimalNumber
          //target: @reportConfig.nps_target
          //targetFormat: noDecimalNumber
          //navigateTo: page_GamingResponses
        }
      }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget dataGrid #dataGridWidget_WinLose {
    label: "Win/Lose by Location"
    size: halfwidth
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "### Did you win or lose during this visit?"

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData

    }


    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_current_counts {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
      //navigateTo: page_RespondentsTable
      //navigateFilter: IN(surveyDataset:NPSVal, "A")
      }

    }

    column #column_NPS {
      label: "NPS®"
      column cut {
        total: none
        value: surveyDataset:WIN_LOSE

        cell #cell {
          value: nps(@reportConfig.nps_qid) * 100
          format: noDecimalNumber
          //extraValue: count(@reportConfig.nps_qid)
          //extraValueFormat: noDecimalNumber
          //target: @reportConfig.nps_target
          //targetFormat: noDecimalNumber
          //navigateTo: page_GamingResponses
        }
      }

    }


    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

  } // end widget
  widget markdown #markdownWidget_6 {
    hide: true
    markdown: "## **Southland Casino Hotel Personas** 
### Based on the question: Why do you visit a regional casino?"

    size: large
  }
  widget dataGrid #dataGridWidget_SouthlandGamingSegmentation {
    label: "Southland Casino Hotel Personas - Why do you visit a regional casino?"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true
    hide: true
    sort rows {
      sortBy: "/Satisfaction_top"
      sortOrder: descending
    }

    row cut {
      value: :GAMING_SEGMENTATION$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:GAMING_SEGMENTATION$value)
        format: noDecimalNumber
        navigateTo: page_SouthlandSegmentationResponses
      }
    }

    column #column_agree {
      label: "% Agree (Top 2)"
      cell {
        value: top2percent(:GAMING_SEGMENTATION$value)
        format: noDecimalPercent
        navigateTo: page_SouthlandSegmentationResponses

      }
    }

    column #AgreePosNegNeutral {
      label: " % Agree Distribution"

      cell microchart {
        value: count(surveyDataset:GAMING_SEGMENTATION$value)
        format: noDecimalNumber

        breakdownBy cut {
          value: recode(:GAMING_SEGMENTATION$value, @sevenPtAgree3cats)
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: noDecimalPercent

        }
      }
    }


    column #column_Agree_Trends {
      label: "Agree Trends (% Top 2)" + " - " + @Gaming_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top2percent(:GAMING_SEGMENTATION$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Gaming_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_SouthlandPersonas {
    label: "Southland Casino Hotel Personas"
    size: halfwidth
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "### Click on any value to see response details"

  //   description: "### Note: To be assigned a persona, all 10 questions had to be answered.

  //  Click on any value to see response details"

    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row cut #row_Southland_segments {
      value: :Southland_Gaming_Seg_assign
      total: none
    }

    column {

      label: "n"


      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        navigateTo: page_SouthlandSegmentationResponses

      }

    }

    column #column_NPS {
      label: "NPS®"

      cell #cell {
        value: nps(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        navigateTo: page_SouthlandSegmentationResponses
      }

    }

    column #column_OSAT {
      label: "OSAT"

      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: noDecimalPercent
        navigateTo: page_SouthlandSegmentationResponses
      }

    }

  } // end widget
} // end page
page #page_KSCVC_Overview {
  label: "Kennedy Space Center"
  //hide: true
  access rules {
    rule claim {
      name: "UserSegment"
      value: "All", "KSCVC"
      //value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_KSCVCSurvey()
    label: "KSCVC survey Only"
  }


  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  // filter expression {
  //   value: _isnull(surveyDataset:hSMGData)
  //   label: "Current Data Only (no historical)"

  // }
  layoutArea toolbar {
    filter multiselect #f_NumVisits {
      label: "Number of Visits"
      optionsFrom: surveyDataset:NO_VISITS
    }
  }
  widget headline #headlineWidget_KSCVC_Overview {

    label: "Voice of Guest Dashboard"

    size: large

    tile markdown #markdownTile_2 {
      value: "# Kennedy Space Center 
### This dashboard compiles Kennedy Space Center survey data collected  via emails sent directly to guests within 1 day post visit. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatim comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a location. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }

    tile button #buttonTile {
      value: "Click here to see information about guest demographics"
      navigateTo: "page_Demos_KSCVC"
      navigateOptions: "same_tab"

      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
    }

  } // end widget
  widget kpi #kpiWidget_Overall_NPS {
    label: "KSCVC NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100

      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_kscvc_target
      //target: parseReal(SitesHierarchySimplified:NPSTarget)
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **Kennedy Space Center Visitors Complex.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "KSCVC OSAT"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_kscvc_target
//target: average(parseReal(SitesHierarchySimplified:OSATTarget), SitesHierarchySimplified:id="1")
    }


    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **Kennedy Space Center Visitors Complex.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  } // end widget
  widget kpi #kpiWidget_Overall_Value {
    label: "KSCVC Value"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top2percent(@reportConfig.value_qid)
      //  value: 35
      label: "Value (Top 2 Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.value_kscvc_target
    }
    infobox #infobox {
      label: "Overall Value"
      info: @reportConfig.value_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.value_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Value KPI for **Kennedy Space Center Visitors Complex.**   The Overall Value KPI is based on the extent to which guests say KSCVC offers an ʺExtremely Goodʺ or ʺVery Goodʺ value. To see more information on Value, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.value_qid))
      label: "Average Value Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.value_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  } // end widget
  widget kpi #kpiWidget_Education {
    label: "Educational Experience at KSCVC"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(:EDUC_EXP.educational)
      //  value: 35
      label: "Educ Exp (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.educ_kscvc_target
    }
    infobox #infobox {
      label: "Education Experience"
      info: "This question assesses the extent to which guests agree that their Kennedy Space Center Visitor Complex offered them an educational experience.

Educational Experience is measured on a five-point scale:

Strongly Disagree
Disagree
Neither Agree Nor Disagree
Agree
Strongly Agree

Where a higher score is better.

We look at value based on the percentage of guests who Strongly Agree."
      size: medium
    }
    tile value #valueTile {
      value: count(:EDUC_EXP.educational)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Educational Experience KPI for **Kennedy Space Center Visitors Complex.**   This metric is based on the extent to which guests ʺStrongly Agreeʺ that KSCVC offered an educational experience. To see more information on this metric, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(:EDUC_EXP.educational))
      label: "Average Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(:EDUC_EXP.educational)
      label: "% Disagree"
      format: percentDefaultFormatter
    }
  } // end widget
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small

    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_11 {
    label: "Recognize a Team Member?"
    hide: true
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  } // end widget
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: primary


      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  } // end widget
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
    }
  } // end widget
  widget headline #headlineWidget_OpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :PROBLEM
    }
    palette: redtogreen2ptscale

    navigateTo: "page_Parks_Overview"
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  } // end widget
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor

    select #KSCVC_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget headline #headlineWidget_KDAs_Location {

    label: "Key Driver Analysis"
    size: large

    select #kscvc_addl_keydrivers_selector {
      label: "Select a Key Driver Analysis"
      options: item {
        label: "Select a Key Driver Analysis"
        value: 0
      },
      item {
        label: "What Drives Satisfaction with KSCVC?"
        value: 1
      },
      item {
        label: "What Drives Attraction Satisfaction?"
        value: 2
      },
      item {
        label: "What Drives Restaurant Satisfaction?"
        value: 3
      },
      item {
        label: "What Drives Premium Experience Satisfaction?"
        value: 4
      },
      item {
        label: "What Drives Gift/Retail Shop Satisfaction?"
        value:5
      }

    }

    tile markdown #markdownTile_2 {
      value: "### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

### There are several analytic views that provide us with strategic direction on what areas to promote as well as those areas that we should consider fixing . To view these, please select  an analysis from the dropdown above."
    }

  } // end widget
  widget keyDrivers #keyDriversWidget_SAT_KSCVC {
    label: "What Drives Satisfaction with KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 1

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: correlation
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis uses correlation to look for patterns in the data to determine how guest experiences influence their overall satisfaction with KSCVC. This shows us where to target improvement in our processes and experiences."
    importanceLimit: 0.3
    dependentVariable: surveyDataset:SAT
    independentVariables: surveyDataset:SAT_EXPERIENCES.attractions, surveyDataset:SAT_EXPERIENCES.bus, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.premiums, surveyDataset:SAT_EXPERIENCES.shops, surveyDataset:SAT_EXPERIENCES.rides
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_KSCVC
  widget keyDrivers #keyDriversWidget_SAT_Attract {
    label: "What Drives Attraction Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 2

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 33
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how experiences with attractions at KSCVC influence their overall attraction satisfaction. This shows us where to target improvement in our attraction processes and experiences."
    importanceLimit: 0.3
    dependentVariable: surveyDataset:SAT_EXPERIENCES.attractions
    independentVariables: surveyDataset:DRILL_ATTRACTION.cleanliness, surveyDataset:DRILL_ATTRACTION.quality, surveyDataset:DRILL_ATTRACTION.staff
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Attract
  widget keyDrivers #keyDriversWidget_SAT_Restaurants {
    label: "What Drives Restaurant Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 3

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 17
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation

      size: large
    }
    description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_EXPERIENCES.restaurants
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.quality, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.staff
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Restaurants
  widget keyDrivers #keyDriversWidget_SAT_Prem_Attract1 {
    label: "What Drives Premium Attraction Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 4

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 33
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with premium attractions influence their overall premium attraction satisfaction. This shows us where to target improvement in our processes and experiences with premium attractions."
    importanceLimit: 0.2
    dependentVariable: surveyDataset:SAT_EXPERIENCES.premiums
    independentVariables: surveyDataset:DRILL_PREMIUM.foodquality, surveyDataset:DRILL_PREMIUM.quality, surveyDataset:DRILL_PREMIUM.staff, surveyDataset:DRILL_PREMIUM.value
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Prem_Attract1
  widget keyDrivers #keyDriversWidget_SAT_Shops1 {
    label: "What Drives Gift/Retail Shop Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 5

    filter expression {
      value: selected(:PURCHASE, "1")

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 25
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the gift/retail shop influence their overall gift/retail shop satisfaction. This shows us where to target improvement in our bar processes and experiences.

### Note: This analysis is for those who indicated they made a purchase."
    importanceLimit: 0.20
    warningText: @reportConfig.kda_warningText
    dependentVariable: surveyDataset:SAT_EXPERIENCES.shops
    independentVariables: surveyDataset:DRILL_SHOPS.value, surveyDataset:DRILL_SHOPS.speed, surveyDataset:DRILL_SHOPS.shopsat, surveyDataset:DRILL_SHOPS.variety, surveyDataset:DRILL_SHOPS.staff, surveyDataset:DRILL_SHOPS.merch
  } // end widget keyDriversWidget_SAT_Shops1
  widget keyDrivers #keyDriversWidget_SAT_Shops2 {
    label: "What Drives Gift/Retail Shop Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 5

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 25
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the gift/retail shop influence their overall gift/retail shop satisfaction. This shows us where to target improvement in our bar processes and experiences.

### Note: This analysis is for those who did not make a purchase."
    importanceLimit: 0.20
    warningText: @reportConfig.kda_warningText
    dependentVariable: surveyDataset:SAT_EXPERIENCES.shops
    independentVariables: surveyDataset:DRILL_SHOPS.shopsat, surveyDataset:DRILL_SHOPS.variety, surveyDataset:DRILL_SHOPS.staff, surveyDataset:DRILL_SHOPS.merch
  } // end widget keyDriversWidget_SAT_Shops2
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  } // end widget
  widget table #tableWidget_comments {
    label: "Visitor Comments"
    size: "large"
    table: surveyDataset:

    showHeader: true
    sortOrder: descending
    sortColumn: comments

    headerNumberOfLines: 3
    stretchColumns: true

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response
    description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response."


    select #OpenEnd_selector {
      label: "Select Question"
      options: item {
        label: "Visit Comments"
        value:  {
          selectQuestion: surveyDataset:VISIT_COMMENTS
          selectFilter: surveyDataset:VISIT_COMMENTS != ""
        }

      },
	    item {
        label: "Restaurant Comments"
        value:  {
          selectQuestion: surveyDataset:RESTAURANT_COMMENTS
          selectFilter: surveyDataset:RESTAURANT_COMMENTS != ""
        }

      },
      item {
        label: "Problem Details"
        value:  {
          selectQuestion: surveyDataset:PROBLEM_DETAIL
          selectFilter: surveyDataset:PROBLEM_DETAIL != ""
        }

      },
      item {
        label: "Team Recognition"
        value:  {
          selectQuestion: surveyDataset:RECOG_DETAIL
          selectFilter: surveyDataset:RECOG_DETAIL != ""
        }

      }    

    } // end OpenEnd_selector
    filter expression {
      value: @OpenEnd_selector.selected.selectFilter
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }


    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }


    column response #comments {
      //sortBy: comment
      //header: "Location: " + surveyDataset:LocationName
      footer: @reportConfig.intvdate
     // width: 300px
      enableColumnFilter: true
      comment: @OpenEnd_selector.selected.selectQuestion

    }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Rec"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    column metric #copy_of_metricColumn {
      label: "OSAT"
      value: score(@reportConfig.osat_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

    column metric #copy_of_metricColumn2 {
      label: "Restaurants Sat"
      value: score(:SAT_EXPERIENCES.restaurants)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

  } // end widget
  widget headline #markdownWidget_PerformanceTrends {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    }

  } // end widget
  widget dataGrid #dataGridWidget_ExperiencesSat {
    label: "Satisfaction with Experiences"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_EXPERIENCES$field
      total: none

    }
    column #column_current_counts {
     // value: count(:SAT_EXPERIENCES$value)
      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:SAT_EXPERIENCES$value)
        navigateTo: "page_KSCVCResponses"
       // showBase: true
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell #undefined {
        format: noDecimalPercent
        value: top1percent(:SAT_EXPERIENCES$value)
        navigateTo: "page_KSCVCResponses"
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_EXPERIENCES$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_AttractionsSat {
    label: "Attractions Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    select #attractions_filter {
      label: "Filter by Attraction Rated"
      mode: multi

      options: @categorySet_attraction_rated.items
    }
    filter expression {
      value: selected(:ATTRACT_INSERT, @attractions_filter.selected)
    }

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_ATTRACTION$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_ATTRACTION$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_ATTRACTION$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_ATTRACTION$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_BusToursSat {
    label: "Bus Tours Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut #Bus {
      value: :DRILL_BUS$field
    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_BUS$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_BUS$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_BUS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RestaurantSat {
    label: "Restaurant Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_RESTAURANT$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_RESTAURANT$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_RESTAURANT$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_PremiumsSat {
    label: "Premium Experience Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    select #premium_exp_filter {
      label: "Filter by Premium Rated"
      mode: multi

      options: @categorySet_premium_exp_rated.items
    }
    filter expression {
      value: selected(:PREMIUM_INSERT, @premium_exp_filter.selected)
    }

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_PREMIUM$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_PREMIUM$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_PREMIUM$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_PREMIUM$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_RetailSat {
    label: "Gift/Retail Shop Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    select #shops_filter {
      label: "Filter by Shop"
      mode: multi

      options: @categorySet_shop_rated.items
    }
    filter expression {
      value: selected(:SHOPS_INSERT, @shops_filter.selected)
    }

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_SHOPS$field
      total: none

    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_SHOPS$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_SHOPS$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_SHOPS$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget headline #headlineWidget_15 {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "# **Guests Experience Profiles**
### These charts show the types of experiences guests reported having while at Kennedy Space Center Visitor Complex. Some of these questions are multi-select and/or are asked of specific sub-segments of guests - these are noted in each chart."
    }

  } //end widget
  widget chart #chartWidget_Tickets {
    label: "Method of Purchasing Tickets"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:TICKETS)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
      textSize: 150
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cut #cutCategory {
      value: :TICKETS
      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "This shows how guests acquired their tickets; each guest was allowed a single answer."
  } //end widget
  widget chart #chartWidget_Reasons {
    label: "Reason for Visit"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:PURPOSE_VISIT)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cut #cutCategory {
      value: :PURPOSE_VISIT
      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "This shows the main reason guests visited Kennedy Space Center Visitor Complex; each guest was allowed a single answer."
  } //end widget
  widget chart #chartWidget_Experiences {
    label: "Guest Experiences During Visit"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:respid)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
      textSize: 225
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cutByMulti #cutCategory {
      value: :EXPERIENCES
      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "This shows the various aspects of Kennedy Space Center Visitor Center that guests experienced during their visit; each guest could pick multiple answers."
    removeEmptyCategories: true
    removeEmptySeries: true
  } //end widget
  widget chart #chartWidget_Attractions {
    label: "Attractions Experienced During Visit"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:respid)
      percentOver: "categories"
      format: percentDefaultFormatter
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cutByMulti #cutCategory {
      value: :ATTRACTIONS_SEEN
      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "Guests randomly selected to evaluate attractions were asked to identify which attractions they visited. Each guest could pick multiple answers."
    removeEmptySeries: true
    removeEmptyCategories: true
  } //end widget
  widget chart #chartWidget_RestaurantsRated {
    label: "Restaurants Rated"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:respid)
      percentOver: "categories"
      format: percentDefaultFormatter
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cut #cutCategory {
      value: :RESTAURANT_INSERT_TEXT
      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "Guests randomly selected to evaluate restaurants were asked to identify which restaurants they visited. Each guest could pick multiple answers."
    removeEmptyCategories: true
    removeEmptySeries: true
  } //end widget
  widget chart #chartWidget_PremiumTours {
    label: "Premium Tours Experienced"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:respid)
      percentOver: "categories"
      format: percentDefaultFormatter
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cutByMulti #cutCategory {
      value: :PREMIUM_PURCHASED

      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "Guests randomly selected to evaluate premium attractions were asked to identify which attractions they visited. Each guest could pick multiple answers."
    removeEmptyCategories: true
    removeEmptySeries: true
  } //end widget
  widget chart #chartWidget_ShopsVisited {
    label: "Gift or Retail Shops Visited"
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:respid)
      percentOver: "categories"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      label: "% of Guests"
      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    category cutByMulti #cutCategory {
      value: :SHOPS_VISITED

      sortOrder: descending
      sortBy: "series"
    }
    size: halfwidth
    description: "Guests randomly selected to evaluate gift and retail shops were asked to identify which locations they visited. Each guest could pick multiple answers."
  } //end widget
  widget dataGrid #dataGridWidget_RestaurantKPIs {
    label: "Restaurant KPIs"
    size: "large"


    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_RatedRestaurant()
      label: "Restaurant Answered"
    }

    row cut {
      value: surveyDataset:RESTAURANT_INSERT_TEXT
      label: "Kennedy Space Center"
  //showLabel: true
      totalLabel: "Kennedy Space Center Visitor Center"
    }

    column #column_restaurant_osat {
      cell #cell {

        value: top1percent(surveyDataset:SAT_EXPERIENCES.restaurants)
        //showBase: true
        format: oneDecimalPercent
        extraValue: count(surveyDataset:SAT_EXPERIENCES.restaurants)
        extraValueFormat: noDecimalNumber

        target: @reportConfig.restaurant_osat_target
        view: comparativeStatisticView
        navigateTo: "page_KSCVCResponses"
      }
      label: "Restaurant OSAT"
    }

    column #column_restaurant_osat_trends {
      cell microchart #cell {
        value: top1percent(surveyDataset:SAT_EXPERIENCES.restaurants)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
        breakdownBy date #dateBreakdownby {
          value: :YieldDateTime
          breakdownBy: @KSCVC_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }
      }
      label: "Restaurant OSAT Trends" + " - " + @KSCVC_Timeframe_Selector.selectedLabel
    }

    column #column_quality {
      label: "Restaurant - Quality"
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.quality)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.quality)
        extraValueFormat: noDecimalNumber
      }
    }
    column #column_value {
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.value)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.value)
        extraValueFormat: noDecimalNumber
      }
      label: "Restaurant - Value"
    }
    column #column_staff {
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.staff)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.staff)
        extraValueFormat: noDecimalNumber
      }
      label: "Restaurant - Staff Friendliness"
    }
    column #column_speed {
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.speed)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.speed)
        extraValueFormat: noDecimalNumber
      }
      label: "Restaurant - Speed"
    }
    column #column_variety {
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.variety)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.variety)
        extraValueFormat: noDecimalNumber
      }
      label: "Restaurant - Variety"
    }
    column #column_clean {
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.cleanliness)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.cleanliness)
        extraValueFormat: noDecimalNumber
      }
      label: "Restaurant - Cleanliness"
    }

    column #column_kiosk {
      cell #cell {
        value: top1percent(surveyDataset:DRILL_RESTAURANT.kiosk)
        format: oneDecimalPercent
        extraValue: count(surveyDataset:DRILL_RESTAURANT.kiosk)
        extraValueFormat: noDecimalNumber
      }
      label: "Restaurant - Kiosk"
    }
    removeEmptyRows: true
    cardTransparent: false
    //description: "Note: Restaurant satisfaction at the individual restaurant level started in June 2023.  The Kennedy Space Center target for Restaurant OSAT is " + @reportConfig.restaurant_osat_target + "%. Satisfaction shown as Top box % based on 5 point scale."
    description: "Note: Restaurant satisfaction at the individual restaurant level started in June 2023.  The Kennedy Space Center goal for Restaurant OSAT is **50%**. Satisfaction shown as Top box % based on 5 point scale."

    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: gridDefaultValueColorFormatter
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }

    showLegend: true
  } //end widget
} // end page
page #page_Lizard_Overview {
  label: "Lizard Island"
  hide: true
  access rules {
    rule claim {
      name: "UserSegment"
      //value: "All", "KSCVC"
      value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_LizardIslandSurvey()
    label: "Lizard Island survey only"
  }


  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  // filter expression {
  //   value: _isnull(surveyDataset:hSMGData)
  //   label: "Current Data Only (no historical)"

  // }
  layoutArea toolbar {
    filter multiselect #f_NumVisits {
      label: "Number of Visits"
      optionsFrom: surveyDataset:NO_VISITS
    }
  }
  widget headline #headlineWidget_KSCVC_Overview {

    label: "Voice of Guest Dashboard"

    size: large

    tile markdown #markdownTile_2 {
      value: "# Lizard Island
### This dashboard compiles Lizard Island survey data collected  via emails sent directly to guests within 1 day post visit. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatim comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a location. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }

    tile button #buttonTile {
      value: "Click here to see information about guest demographics"
      navigateTo: "page_Demos_LizardIsland"
      navigateOptions: "same_tab"

      navigateFilter: surveyDataset:filterMeasure_LizardIslandSurvey()
    }

  } // end widget
  widget kpi #kpiWidget_Overall_NPS {
    label: "Lizard Island NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100

      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_kscvc_target
      //target: parseReal(SitesHierarchySimplified:NPSTarget)
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **Lizard Island.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Lizard Island OSAT"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_kscvc_target
//target: average(parseReal(SitesHierarchySimplified:OSATTarget), SitesHierarchySimplified:id="1")
    }


    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **Lizard Island.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  } // end widget
  widget kpi #kpiWidget_Overall_Value {
    label: "Lizard Island Value"
    size: small

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top2percent(@reportConfig.value_qid)
      //  value: 35
      label: "Value (Top 2 Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.value_kscvc_target
    }
    infobox #infobox {
      label: "Overall Value"
      info: @reportConfig.value_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.value_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Value KPI for **Lizard Island.**   The Overall Value KPI is based on the extent to which guests say KSCVC offers an ʺExtremely Goodʺ or ʺVery Goodʺ value. To see more information on Value, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.value_qid))
      label: "Average Value Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.value_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  } // end widget
  widget headline #headlineWidget_Problem {
    label: "Problem During Visit?"
    hide: true
    size: small

    tile text #textTile {
      value: "1) % Visitors That Indicated a Problem During Visit:"
      fontSize: 20
    }

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1") / count(surveyDataset:) * 100
      valueFormatter: noDecimalPercent

      //valueColorFormatter: gaugeDefaultColorFormatter_V2
      fontSize: 35
    }
    tile value #valueTile__base {
      value: count(surveyDataset:, surveyDataset:PROBLEM = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_2 {
      value: "2) % Visitors That Reported a Problem During Visit:"
      fontSize: 20
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1") / count(surveyDataset:) * 100
      fontSize: 35
      valueFormatter: noDecimalPercent
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_3__base {
      value: count(surveyDataset:, surveyDataset:PROB_REPORTED = "1")
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile text #textTile_3 {
      value: "3)  Satisfaction (% Top Box) with Problem Resolution:"
      fontSize: 20
    }

    tile value #valueTile_4 {
      value: top1percent(:RESOLUTION_SAT)
      fontSize: 35
      valueFormatter: percentDefaultFormatter
      //valueColorFormatter: gaugeDefaultColorFormatter_V2
    }
    tile value #valueTile_4__base {
      value: count(:RESOLUTION_SAT)
      pretext: "Responses: "
      fontSize: 14
      spacing: "none"
      valueFormatter: noDecimalNumber
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_ProblemDrilldown"
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
      type: danger
      navigateOptions: "same_tab"
    }


    infobox #infobox {
      label: ""
      info: ""
    }
  } // end widget
  widget headline #headlineWidget_11 {
    label: "Recognize a Team Member?"
    hide: true
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors recognized a Team Member"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1") / count(surveyDataset:TEAM_REC) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }

    tile button #buttonTile {
      value: "Learn More"
      navigateTo: page_TeamRecog
      navigateFilter: IN(surveyDataset:PROBLEM, "1") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: primary
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:TEAM_REC = "1")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  } // end widget
  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: primary


      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_KSCVCSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  } // end widget
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
    }
  } // end widget
  widget headline #headlineWidget_OpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :PROBLEM
    }
    palette: redtogreen2ptscale

    navigateTo: "page_Parks_Overview"
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  } // end widget
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_KSCVCSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor

    select #Lizard_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Lizard_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent
        //showBase: true
        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal

      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Lizard_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Lizard_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Lizard_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
//   widget headline #headlineWidget_KDAs_Location {

//     label: "Key Driver Analysis"
//     size: large

//     select #lizard_addl_keydrivers_selector {
//       label: "Select a Key Driver Analysis"
//       options: item {
//         label: "Select a Key Driver Analysis"
//         value: 0
//       },
//       item {
//         label: "What Drives Satisfaction with Lizard Island?"
//         value: 1
//       }
//       // item {
//       //   label: "What Drives Attraction Satisfaction?"
//       //   value: 2
//       // },
//       // item {
//       //   label: "What Drives Restaurant Satisfaction?"
//       //   value: 3
//       // },
//       // item {
//       //   label: "What Drives Premium Experience Satisfaction?"
//       //   value: 4
//       // },
//       // item {
//       //   label: "What Drives Gift/Retail Shop Satisfaction?"
//       //   value:5
//       // }

//     }

//     tile markdown #markdownTile_2 {
//       value: "### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

// ### There are several analytic views that provide us with strategic direction on what areas to promote as well as those areas that we should consider fixing . To view these, please select  an analysis from the dropdown above."
//     }

//   } // end widget
  widget keyDrivers #keyDriversWidget_SAT_LizardIsland {
    label: "What Drives Satisfaction with Lizard Island?"
    //hide: @lizard_addl_keydrivers_selector.selected != 1
    hide: true
    //minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    minimumSampleSize: 1
    algorithm: correlation
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_correlation
      info: @reportConfig.kda_infobox_info_correlation

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis uses correlation to look for patterns in the data to determine how guest experiences influence their overall satisfaction with KSCVC. This shows us where to target improvement in our processes and experiences."
    importanceLimit: 0.3
    dependentVariable: surveyDataset:SAT
    independentVariables: surveyDataset:SAT_RESORT_EXPERIENCES_transfer, surveyDataset:SAT_RESORT_EXPERIENCES_aquatic_tours, surveyDataset:SAT_RESORT_EXPERIENCES_aquatic_activities, surveyDataset:SAT_RESORT_EXPERIENCES_spa, surveyDataset:SAT_RESORT_EXPERIENCES_athletic, surveyDataset:SAT_RESORT_EXPERIENCES_nature, surveyDataset:SAT_RESORT_EXPERIENCES_scuba
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_KSCVC
  widget keyDrivers #keyDriversWidget_SAT_Attract {
    label: "What Drives Attraction Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 2

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 33
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how experiences with attractions at KSCVC influence their overall attraction satisfaction. This shows us where to target improvement in our attraction processes and experiences."
    importanceLimit: 0.3
    dependentVariable: surveyDataset:SAT_EXPERIENCES.attractions
    independentVariables: surveyDataset:DRILL_ATTRACTION.cleanliness, surveyDataset:DRILL_ATTRACTION.quality, surveyDataset:DRILL_ATTRACTION.staff
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Attract
  widget keyDrivers #keyDriversWidget_SAT_Restaurants {
    label: "What Drives Restaurant Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 3

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 17
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation

      size: large
    }
    description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_EXPERIENCES.restaurants
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.quality, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.staff
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Restaurants
  widget keyDrivers #keyDriversWidget_SAT_Prem_Attract1 {
    label: "What Drives Premium Attraction Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 4

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 33
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with premium attractions influence their overall premium attraction satisfaction. This shows us where to target improvement in our processes and experiences with premium attractions."
    importanceLimit: 0.2
    dependentVariable: surveyDataset:SAT_EXPERIENCES.premiums
    independentVariables: surveyDataset:DRILL_PREMIUM.foodquality, surveyDataset:DRILL_PREMIUM.quality, surveyDataset:DRILL_PREMIUM.staff, surveyDataset:DRILL_PREMIUM.value
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Prem_Attract1
  widget keyDrivers #keyDriversWidget_SAT_Shops1 {
    label: "What Drives Gift/Retail Shop Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 5

    filter expression {
      value: selected(:PURCHASE, "1")

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 25
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the gift/retail shop influence their overall gift/retail shop satisfaction. This shows us where to target improvement in our bar processes and experiences.

### Note: This analysis is for those who indicated they made a purchase."
    importanceLimit: 0.20
    warningText: @reportConfig.kda_warningText
    dependentVariable: surveyDataset:SAT_EXPERIENCES.shops
    independentVariables: surveyDataset:DRILL_SHOPS.value, surveyDataset:DRILL_SHOPS.speed, surveyDataset:DRILL_SHOPS.shopsat, surveyDataset:DRILL_SHOPS.variety, surveyDataset:DRILL_SHOPS.staff, surveyDataset:DRILL_SHOPS.merch
  } // end widget keyDriversWidget_SAT_Shops1
  widget keyDrivers #keyDriversWidget_SAT_Shops2 {
    label: "What Drives Gift/Retail Shop Satisfaction at KSCVC?"
    hide: @kscvc_addl_keydrivers_selector.selected != 5

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: 25
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 90
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: halfwidth
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the gift/retail shop influence their overall gift/retail shop satisfaction. This shows us where to target improvement in our bar processes and experiences.

### Note: This analysis is for those who did not make a purchase."
    importanceLimit: 0.20
    warningText: @reportConfig.kda_warningText
    dependentVariable: surveyDataset:SAT_EXPERIENCES.shops
    independentVariables: surveyDataset:DRILL_SHOPS.shopsat, surveyDataset:DRILL_SHOPS.variety, surveyDataset:DRILL_SHOPS.staff, surveyDataset:DRILL_SHOPS.merch
  } // end widget keyDriversWidget_SAT_Shops2
  widget headline #headlineWidget_Comments {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  } // end widget
  widget table #tableWidget_comments {
    label: "Visitor Comments"
    size: "large"
    table: surveyDataset:

    showHeader: true
    sortOrder: descending
    sortColumn: comments

    headerNumberOfLines: 3
    stretchColumns: true

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response
    description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response."


    select #OpenEnd_selector {
      label: "Select Question"
      options: item {
        label: "Visit Comments"
        value:  {
          selectQuestion: surveyDataset:VISIT_COMMENTS
          selectFilter: surveyDataset:VISIT_COMMENTS != ""
        }

      },
      	    item {
        label: "Lodging Comments"
        value:  {
          selectQuestion: surveyDataset:LODGING_COMMENTS
          selectFilter: surveyDataset:LODGING_COMMENTS != ""
        }

      },
	    item {
        label: "Restaurant Comments"
        value:  {
          selectQuestion: surveyDataset:RESTAURANT_COMMENTS
          selectFilter: surveyDataset:RESTAURANT_COMMENTS != ""
        }

      },
      	    item {
        label: "Experiences Comments"
        value:  {
          selectQuestion: surveyDataset:EXPERIENCES_COMMENTS
          selectFilter: surveyDataset:EXPERIENCES_COMMENTS != ""
        }

      },
      item {
        label: "Problem Details"
        value:  {
          selectQuestion: surveyDataset:PROBLEM_DETAIL
          selectFilter: surveyDataset:PROBLEM_DETAIL != ""
        }

      },
      item {
        label: "Team Recognition"
        value:  {
          selectQuestion: surveyDataset:RECOG_DETAIL
          selectFilter: surveyDataset:RECOG_DETAIL != ""
        }

      }    

    } // end OpenEnd_selector
    filter expression {
      value: @OpenEnd_selector.selected.selectFilter
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }


    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }


    column response #comments {
      //sortBy: comment
      header: "Location: " + surveyDataset:LocationName
      footer: @reportConfig.intvdate
     // width: 300px
      enableColumnFilter: true
      comment: @OpenEnd_selector.selected.selectQuestion

    }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Rec"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    column metric #copy_of_metricColumn {
      label: "OSAT"
      value: score(@reportConfig.osat_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

    column metric #copy_of_metricColumn2 {
      label: "Restaurants Sat"
      value: score(:DRILL_RESTAURANT.restaurant)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

  } // end widget
  widget headline #markdownWidget_PerformanceTrends {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    }

  } // end widget
  widget dataGrid #dataGridWidget_ExperiencesSat {
    label: "Satisfaction with Experiences"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_RESORT_EXPERIENCES$field
      total: none

    }
    column #column_current_counts {

      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:SAT_RESORT_EXPERIENCES$value)
        navigateTo: "page_KSCVCResponses"
       // showBase: true
      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell #undefined {
        format: noDecimalPercent
        value: top1percent(:SAT_RESORT_EXPERIENCES$value)
        navigateTo: "page_KSCVCResponses"
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lizard_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_RESORT_EXPERIENCES$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lizard_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_LodgingSat {
    label: "Lodging Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut #Lodging {
      value: :DRILL_LODGING$field
      total: none
    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_LODGING$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lizard_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lizard_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RoomSat {
    label: "Room Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut #Lodging {
      value: :DRILL_ROOM$field
      total: none
    }
    column #column_current_counts {
      label: "Number of Responses"
      cell {
        value: count(:DRILL_ROOM$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lizard_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lizard_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RestaurantSat {
    label: "Restaurant Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_RESTAURANT$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_RESTAURANT$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_RESTAURANT$value)
        format: noDecimalNumber
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        navigateTo: "page_KSCVCResponses"

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Lizard_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Lizard_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }

    }

  } //end widget
} // end page
page #page_AustraliaOverview {
  label: "Australia Locations"
  hide: true
  access rules {
    rule claim {
      name: "UserSegment"
      //value: "All", "Lodging", "Parks"
      value: "Test"
    }
  }

  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_AustraliaLocations()
    label: "Australia Page Locations"
  }


  filter expression #NPSAnswered2 {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }


  widget headline #headlineWidget_Lodging_Overview {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Australia Overview 
### This dashboard compiles lodging survey data collected  via emails sent directly to guests within 1 day post visit. 
 
Included in the report is a view of: 
- Key performance indicators: NPS® and Overall Satisfaction 
- Key drivers of satisfaction
- Trends
- Verbatim comments from guests
 
You can click on the filter icon in the upper left-hand corner of the report to refine your dashboard, including narrowing your focus to a location. When filtering results, please exercise caution in interpretation of scores when the number of records is below 50.

***By default, this report looks at only the current year to date; to review trend data prior to the current year, please remove this filter (or customize the filter to a time range of your choosing). Goals and targets are based on current year targets.***"

    }

    tile text #textTile {
      value: "Your assigned location(s):"
      fontSize: 20

    }
    tile value #valueTile_ReportBase {
      filter expression {
        value: _isNull(FromAncestor(SitesHierarchy:^hierarchy, SitesHierarchy:id))
      }
      value: AggText(SitesHierarchy:language_text, ", ", SitesHierarchy:__row_order)
      fontSize: 25

    }

    tile button #buttonTile {
      value: "Click here to see information about guest demographics"
      navigateTo: "page_Demos"
      navigateOptions: "same_tab"

      navigateFilter: surveyDataset:filterMeasure_AustraliaLocations()
    }
    label: "Voice of Guest Dashboard"
  }
  widget kpi #kpiWidget_Overall_NPS {
    label: "Overall Subsidiary NPS®"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }
    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
     // target: @reportConfig.nps_lodging_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **All Australia lodging locations within Parks & Resorts.**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Overall_OSAT {
    label: "Overall Subsidiary OSAT"
    size: small
    ignoreFilters: f_Location

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      target: @reportConfig.osat_lodging_target
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **All Australia lodging locations within Parks & Resorts.**   The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }
  widget kpi #kpiWidget_Location_NPS {
    label: "My Location(s) NPS®"
    size: small

    tile kpi #kpiTile {
      value: nps(@reportConfig.nps_qid) * 100
      //  value: 35
      label: "NPS"

      format: noDecimalNumber
      min: -100
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
      //target: @reportConfig.nps_travel_target
    }
    infobox #infobox {
      label: "NPS®"
      info: @reportConfig.nps_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.nps_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Net Promoter Score® for **your specific Australian Parks & Resorts location(s).**  The Net Promoter Score® is based on the extent to which guests agree that they would recommend us based on a 0-10 scale, where 0 = Not At All Likely and 10 = Extremely Likely. To see more information on NPS®, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:NPS))
      label: "Average Recommendation Score"
      min: 0
      max: 10
      format: twoDecimalNumber
    }
  }
  widget kpi #kpiWidget_Location_OSAT {
    label: "My Location(s) OSAT"
    size: small


    tile kpi #kpiTile {
      value: top1percent(@reportConfig.osat_qid)
      //  value: 35
      label: "OSAT (Top Box)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
       //target: @reportConfig.osat_travel_target     
    }
    infobox #infobox {
      label: "Overall Satisfaction"
      info: @reportConfig.osat_infoText
      size: medium
    }
    tile value #valueTile {
      value: count(@reportConfig.osat_qid)
      label: "Responses"
      format: noDecimalNumber
    }
    description: "This shows our Overall Satisfaction KPI for **your specific Australian Parks & Resorts location(s).**  The Overall Satisfaction KPI is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above.
"
    tile value #valueTile_2 {
      value: average(numeric(@reportConfig.osat_qid))
      label: "Average Satisfaction Score"
      min: 0
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(@reportConfig.osat_qid)
      label: "% Dissatisfied"
      format: percentDefaultFormatter
    }
  }



  widget headline #headlineWidget_NPS_Cats {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Breakdown of Net Promoter Categories**
### The Net Promoter Score, or NPS®, is a metric that describes how likely guests are to recommend us to friends and family. It is seen as a leading indicator of future financial success."
    }

  }

  widget headline #headlineWidget_activePromoters {
    label: "Active Promoters"
    size: small
    //navigateTo: ResponsesModel

    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }

    tile text #textTile {
      value: "of our visitors are Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
      view: iconView
      colorFormatter: NPS_promoters
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_promoters
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "A") AND surveyDataset:filterMeasure_LodgingSurvey()
      type: primary


      navigateOptions: "same_tab"
    }

    view numeric #numericView_infographicTile {
      max: 100
    }

    tile text #textTile_3 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_3 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "A")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }

  } // end widget
  widget headline #headlineWidget_Passives {
    label: "Passives"
    size: small
   // navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "B") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_passives
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "B") AND surveyDataset:filterMeasure_LodgingSurvey()
      type: success
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      fontSize: 24
      valueFormatter: noDecimalNumber
      value: count(surveyDataset:, surveyDataset:NPSVal = "B")
    }
  } // end widget
  widget headline #headlineWidget_Detractors {
    label: "Detractors"
    size: small
    //navigateTo: ResponsesModel
    tile value #valueTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      valueFormatter: noDecimalPercent
    }
    tile text #textTile {
      value: "of our visitors are Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C") / count(surveyDataset:NPSVal) * 100
      view: "iconView_infographicTile"
      colorFormatter: NPS_detractors
    }

    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "horizontal"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    tile button #buttonTile {
      value: "Learn More"
      navigateTo: "page_NPSResponses"
      navigateFilter: IN(surveyDataset:NPSVal, "C") AND surveyDataset:filterMeasure_LodgingSurvey()
      type: danger
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Responses"
      fontSize: 16
    }
    tile value #valueTile_2 {
      value: count(surveyDataset:, surveyDataset:NPSVal = "C")
      fontSize: 24
      valueFormatter: noDecimalNumber
    }
  } // end widget
  widget markdown #markdownWidget_NPS_descrip {
    markdown: "### **NPS® description**
Based on your recent visit, how likely are you to recommend [Location] to a friend or family member?
![NPS description](https://cdn.us.confirmit.com/isa/LDEBDRJXGRLRIIIBIYJTMYHPHPMVLANH/NPS%20visual.png)"
  }
  widget headline #headlineWidget_AM_descript {
    size: small

    tile markdown #markdownTile_2 {
      value: "## **Summary of Action Management Cases**
### We have action cases that are triggered based on guest feedback. This section of the dashboard summarizes the cases that have been created.  "

    }
    tile button #buttonTile {
      value: "Go To Action Management"
      navigateTo: "page_CasesOverview"
      navigateOptions: "same_tab"
      navigateFilter: surveyDataset:filterMeasure_AustraliaLocations()
    }
  }
  widget headline #headlineWidget_totalOpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_InProgressCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #headlineWidget_OverdueCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #chartWidget_Problem {
    label: "Problem During Visit?"
    //hide: true
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      navigateTo: page_ProblemDrilldown
      navigateFilter: surveyDataset:filterMeasure_AustraliaLocations()
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :PROBLEM
    }
    palette: redtogreen2ptscale

   // navigateTo: "page_Parks_Overview"
    description: "To see more details (like who has requested contact and other useful information), please click the appropriate slice of the pie."
  }
  widget chart #chartWidget_TeamRecog {
    label: "Recognize a Team Member?"
    //hide: true
    series #series {
      value: count(:TEAM_REC)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      navigateTo: page_TeamRecog
      navigateFilter: surveyDataset:filterMeasure_AustraliaLocations()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"
    category cut #cutCategory {
      value: :TEAM_REC
    }

    palette: copy_of_greentored2ptscale
    description: "To see guest feedback on team members, please click in the green slice of the pie (the ʺYes, want to recognizeʺ slice)."
  }
  widget headline #headlineWidget_TrendSelector {
    label: "Trends"
    size: large
    cardBackground: @reportConfig.selector_CardBackgroundColor


    select #Australia_Timeframe_Selector {
      label: "Select Timeframe"

      options: @valueSet_date_ranges_1.items

    } // end selector
    tile markdown #markdownTile {
      value: "### Use this selector to see trends in various timeframes"
    }


  }
  widget chart #chartWidget_NPS_Trends_Bars {
    label: "NPS® Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
   // ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @NPS_Timeframe_Selector2.selected.selectFilter
    // }

    // select #NPS_Timeframe_Selector2 {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series_npsCategories {

      value: count(@reportConfig.nps_qid)
      isSecondary: true
      format: noDecimalNumber
      palette: nps_palette_reversed
      chart bar {
        mode: stacked100Percent
        dataLabel: percent

        maxBarSize: 50
        showValue: true

      }
      breakdownBy cut {
        value: :NPSVal
      }

      label: "NPS® Categories"
    }

    series #series_nps {

      value: nps(@reportConfig.nps_qid) * 100
      isSecondary: false
      format: noDecimalNumber
      palette: nps_and_cats_palette
      chart line #lineChart {
        dotSize: 5
        lineWidth: 3
        dotColorFormat: dotColorFormatter
        showDotValue: true

      }
      label: "NPS®"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter

    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100

    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Bars {
    label: "OSAT Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
    // label: @Tkpiselect.selected.kpiLabel + " Trends"   
    palette: kpi_palette
    //ignoreFilters: reportingPeriodFilter

    // filter expression {
    //   value: @OSAT_Timeframe_Selector2.selected.selectFilter
    // }

    // select #OSAT_Timeframe_Selector2 {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items
    // } // end selector
    series #series_osat {
      chart bar #barChart {
        //showBase: true
        maxBarSize: 50
      }
      value: top1percent(@reportConfig.osat_qid)
      isSecondary: false
      format: oneDecimalPercent
      label: "Overall Satisfaction"
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalPercent
      label: "Top Box % (5's)"

      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "Top 2 Box % "
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 60
    }

    base #base {
      value: count(@reportConfig.osat_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
    description: "Note: When sample size is under 50, please review with caution."
  } // end widget
  widget dataGrid #dataGridWidget_LocationKPIs {
    label: "Location KPIs"
    size: large
    ignoreFilters: f_Location
    removeEmptyRows: true
    description: "This view displays a breakdown of the performance of all locations on our key performance indicators. This provides insight on how locations perform in a relative context.
#### **Goals shown are current year goals; please keep this in mind if you change the reporting period.**
"

    filter expression {
      value: count(:, selected(:survey_pid, @reportConfig.surveypid_lizard), SitesHierarchySimplified:^hierarchy) > 0 OR count(:, selected(:survey_pid, @reportConfig.surveypid_gaming), SitesHierarchySimplified:^hierarchy) > 0 OR count(:, selected(:survey_pid, @reportConfig.surveypid_lodging), SitesHierarchySimplified:^hierarchy) > 0

    }

    view comparativeStatistic #view_diff_goal {
      backgroundColorFormatter: background_diff_goal
      valueColorFormatter: text_diff_goal
    }

    row comparison #comparisonRow {
      reportingHierarchy: SitesHierarchySimplified
      showTotal: false
    }

    column #column_current_counts {

      label: "n"

      cell {
        value: count(@reportConfig.nps_qid)
        format: noDecimalNumber
        //navigateTo: page_LodgingResponses

      }

    }

    column #column_current_NPS {

      label: "NPS®"

      // scope reportingPeriod {
      //   period: Current
      // }
      cell {
        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber

        //navigateTo: page_LodgingResponses
       // view: comparativeStatisticView
      }
    }

    column cut #column_Promoters {
      //value: recode(@reportConfig.nps_qid, @NPScats)
      value: surveyDataset:NPSVal
      categories: "'A'"
      label: "Promoters"
      total: none
      cell columnPercentage {
        value: count(@reportConfig.nps_qid)
        format: oneDecimalPercent
       // target: @reportConfig.promoters_target
        extraValue: count(@reportConfig.nps_qid)
        extraValueFormat: noDecimalNumber
        //navigateTo: page_LodgingResponses
        //navigateFilter: IN(surveyDataset:NPSVal, "A")

      }
    }

    column #NPSPosNegNeutral {
      label: " % within NPS® category "

      cell microchart {
        value: count(surveyDataset:)
        format: noDecimalNumber
              //extraValue: count(@reportConfig.nps_qid)
        breakdownBy cut {
          value: surveyDataset:NPSVal

         // value: LoyaltyGrid:value
        }
        microchart stacked100PercentBar {
          valuePosition: none
          palette: nps_palette_reversed
          notAnswered: false
          showTooltip: true
          percentFormat: oneDecimalPercent

        }
      }
    }

    column #column_NPS_Trends {
      label: "NPS® Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
      // filter expression {
      //   value: @Lodging_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart {

        value: NPS(@reportConfig.nps_qid) * 100
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
          //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA


        }
      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }
    }



    column #column_current_OSAT {
      cell #cell {
        value: top1percent(@reportConfig.osat_qid)
        //target: @reportConfig.osat_target
        format: oneDecimalPercent
        showBase: true
        //navigateTo: page_LodgingResponses
        //navigateFilter: _isnotnull(@reportConfig.osat_qid)
      }
      label: "Overall Sat"
    }

    column #column_OSATGoal {

      label: "OSAT Goal"

      format: noDecimalNumber

      cell {

        value: parseReal(SitesHierarchySimplified:OSATTarget)
        format: noDecimalNumber

        //view: comparativeStatisticView
      }
    }


    column #column_OSAT_diff {

      value: surveyDataset:
      total: none

      cell diff {

        main: column_current_OSAT
        other: column_OSATGoal
        diff: absolute
        format: noDecimalNumber
        view: view_diff_goal
      }

      label: "vs. Goal"

    }

    column #column_OSAT_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      // filter expression {
      //   value: @Lodging_Timeframe_Selector.selected.selectFilter
      // }

      cell microchart #cell {
        value: top1percent(@reportConfig.osat_qid)
        format: oneDecimalPercent
        useOnlyExistingColumns: true
        microchart line #barMicrochart {
          min: auto
          max: auto
        }
        breakdownBy date #dateBreakdownby {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        }

      }
      // scope reportingPeriod #reportingPeriodScope {
      //   period: "allData"
      // }

    }

    infobox #infobox {
      label: "Sites KPIs info"
      info: "Color formatting based on target values for the associated KPI. "
    }
    showLegend: true
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }


  } // end widget
  widget headline #headlineWidget_KDAs_Location {
    label: "Key Driver Analysis By Location"
    size: large
    hide: true
    tile markdown #markdown1 {
      value: "### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

### The data below show the relationships at high levels as well as at functional levels."

//### **Please note:** These analyses require a minimum of 100 records to run; if less than 100 records are available, the report will generate an error message. If you see the message 'The accuracy of the model shown falls below the criteria specified. Please exercise caution in the use of these data.' this means that the R-squared value of the model falls below 0.5."

    }

    select #Australian_Locations_Selector {
      label: "Select a Australian Location"

      options: @valueSet_australia_locations.items

    } // end selector
  }
//   widget markdown #markdownWidget_3 {
//     markdown: "## **Key Driver Analysis**

// ### **Key Driver Analysis** provides insight into what influences guests' ratings on our KPIs. Understanding these relationships, combined with an assessment of our performance, provides strategic insights on where we should focus improvement efforts and strengths to promote.

// ### The data below show the relationships at high levels as well as at functional levels. "
//     size: large
//   }

  // widget keyDrivers #keyDriversWidget_NPS_Lodging_Overall {
  //   label: "What Drives Likelihood to Recommend for Lodging Overall?"

  // //attributes removed for this KDA: none
  // //this kda applies to lodging as a whole

  //   hide: @Lodging_Locations_Selector.selected != "Lodging"
  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

  //   minimumSampleSize: @reportConfig.KDAMinimumSampleSize
  //   algorithm: correlation
  //   satisfactionLimit: 80
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: @reportConfig.kda_descriptionText
  //   importanceLimit: 0.5
  //   dependentVariable: surveyDataset:NPS
  //   independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.concierge, surveyDataset:SAT_EXPERIENCES.otheramenities, surveyDataset:SAT_EXPERIENCES.spa, surveyDataset:SAT_EXPERIENCES.shops

  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_NPS_Lodging_Overall

  widget keyDrivers #keyDriversWidget_NPS_Lodging1 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

  //attributes removed for this KDA: breakfast
  //this kda applies to following locations:
    //474A	The Lodge at Tenaya 
    //474B	The Cottages at Tenaya
    //474C	The Explorer Cabins at Tenaya  

    hide: @Lodging_Locations_Selector.selected != "474A" AND @Lodging_Locations_Selector.selected != "474B" AND @Lodging_Locations_Selector.selected != "474C"
    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.concierge, surveyDataset:SAT_EXPERIENCES.otheramenities, surveyDataset:SAT_EXPERIENCES.spa, surveyDataset:SAT_EXPERIENCES.shops

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging1
  widget keyDrivers #keyDriversWidget_NPS_Lodging2 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, spa, other amenities
   //this kda applies to following locations:
    //59841	Peaks of Otter
    //59989A	John Muir Lodge - Kings Canyon National Park
    //59989B	Grant Grove Cabins - Kings Canyon National Park
    //63108	Yavapai Lodge - Grand Canyon National Park
    //63275	Trailer Village RV Park - Grand Canyon National Park

    hide: @Lodging_Locations_Selector.selected != "59841" AND @Lodging_Locations_Selector.selected != "59989A" AND @Lodging_Locations_Selector.selected != "59989B" AND @Lodging_Locations_Selector.selected != "63108" AND @Lodging_Locations_Selector.selected != "63275"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.shops

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging2
  widget keyDrivers #keyDriversWidget_NPS_Lodging3 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, spa
   //this kda applies to following locations:
    //22005A	The Lodge at Geneva on the Lake
    //22005B	The Cottages at Geneva on the Lake
    //58866	Big Meadows Lodge - Shenandoah
    //58867	Skyland Resort - Shenandoah

    hide: @Lodging_Locations_Selector.selected != "22005A" AND @Lodging_Locations_Selector.selected != "22005B" AND @Lodging_Locations_Selector.selected != "58866" AND @Lodging_Locations_Selector.selected != "58867"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.shops, surveyDataset:SAT_EXPERIENCES.otheramenities

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging3
  widget keyDrivers #keyDriversWidget_NPS_Lodging4 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, spa, bars, other amenities
   //this kda applies to following locations:
    //404	Wuksachi Lodge - Sequoia National Park   
    //58148	Kalaloch Lodge
    //59988	Cedar Grove Lodge - Kings Canyon National Park

    hide: @Lodging_Locations_Selector.selected != "404" AND @Lodging_Locations_Selector.selected != "58148" AND @Lodging_Locations_Selector.selected != "59988"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.shops

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging4
  widget keyDrivers #keyDriversWidget_NPS_Lodging5 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, bars, other amenities
   //this kda applies to following locations:
    //139	The Gideon Putnam

    hide: @Lodging_Locations_Selector.selected != "139"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.shops, surveyDataset:SAT_EXPERIENCES.spa

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging5
  widget keyDrivers #keyDriversWidget_NPS_Lodging6 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: concierge, restaurants, bars, shops, spa
   //this kda applies to following locations:
    //28577	Gray Wolf Inn & Suites
    //28578	Yellowstone Park Hotel


    hide: @Lodging_Locations_Selector.selected != "28577" AND @Lodging_Locations_Selector.selected != "28578"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.breakfast, surveyDataset:SAT_EXPERIENCES.otheramenities

    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_NPS_Lodging6
  widget keyDrivers #keyDriversWidget_NPS_Lodging7 {
    label: "What Drives Likelihood to Recommend at " + @Lodging_Locations_Selector.selectedLabel + "?"

   //attributes removed for this KDA: breakfast, concierge, restaurants, bars, shops, spa
   //this kda applies to following locations:
    //59396	The Explorer Cabins at Yellowstone

    hide: @Lodging_Locations_Selector.selected != "59396"

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)
    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: @reportConfig.kda_descriptionText
    importanceLimit: 0.5
    dependentVariable: surveyDataset:NPS
    independentVariables: surveyDataset:Value, surveyDataset:SAT_EXPERIENCES.lodging, surveyDataset:SAT_EXPERIENCES.otheramenities

    warningText: @reportConfig.kda_warningText
    //rSquaredLimit: 0.5
  } // end widget keyDriversWidget_NPS_Lodging7
  widget headline #headlineWidget_KDAs_Location_Addtl {

    label: "Additional Key Driver Analyses for " + @Lodging_Locations_Selector.selectedLabel + ""
    size: large
    hide: true

    select #lodging_addl_keydrivers_selector {
      label: "Select an Additional Key Driver Analysis"
      options: item {
        label: "Select to see other Key Driver Analyses"
        value: 0
      },
      item {
        label: "What Drives Satisfaction with Lodging?"
        value: 1
      },
      item {
        label: "How Do Room Features Impact Lodging Satisfaction?"
        value: 2
      },
      item {
        label: "What Drives Restaurant Satisfaction?"
        value: 3
      },
      item {
        label: "What Drives Bar Satisfaction?"
        value: 4
      }

    }

    tile markdown #markdownTile_2 {
      value: "### There are several analytic views that provide us with strategic direction on what areas to promote as well as those areas that we should consider fixing . To view these, please select  an analysis from the dropdown above."
    }

  }

  // widget keyDrivers #keyDriversWidget_SAT_Lodging_Overall {
  //   label: "What Drives Satisfaction with Lodging Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 1 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

  //   minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    // algorithm: regression
    //// algorithm: correlation

  //   satisfactionLimit: 85
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
  //   importanceLimit: 0.15
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
  //   independentVariables: surveyDataset:DRILL_LODGING.accuracy, surveyDataset:DRILL_LODGING.arrival, surveyDataset:DRILL_LODGING.avail, surveyDataset:DRILL_LODGING.cleanliness, surveyDataset:DRILL_LODGING.staff, surveyDataset:DRILL_LODGING.departure, surveyDataset:DRILL_LODGING.service
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Lodging_Overall

  widget keyDrivers #keyDriversWidget_SAT_Lodging {
    label: "What Drives Satisfaction with Lodging at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 1

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how guest experiences influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
    independentVariables: surveyDataset:DRILL_LODGING.accuracy, surveyDataset:DRILL_LODGING.arrival, surveyDataset:DRILL_LODGING.avail, surveyDataset:DRILL_LODGING.cleanliness, surveyDataset:DRILL_LODGING.staff, surveyDataset:DRILL_LODGING.departure, surveyDataset:DRILL_LODGING.service
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Lodging
  // widget keyDrivers #keyDriversWidget_SAT_Room_Overall {
  //   label: "How Do Room Features Impact Lodging Satisfaction Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 2 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

    // algorithm: regression
    //// algorithm: correlation
  //   satisfactionLimit: 85
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how room features, experiences and characteristics influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
  //   importanceLimit: 0.10
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
  //   independentVariables: surveyDataset:DRILL_ROOM.ac, surveyDataset:DRILL_ROOM.bathamenities, surveyDataset:DRILL_ROOM.bathclean, surveyDataset:DRILL_ROOM.bathfeatures, surveyDataset:DRILL_ROOM.bed, surveyDataset:DRILL_ROOM.cleanliness, surveyDataset:DRILL_ROOM.furnishings, surveyDataset:DRILL_ROOM.quiet, surveyDataset:DRILL_ROOM.smell, surveyDataset:DRILL_ROOM.wifi
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Room_Overall

  widget keyDrivers #keyDriversWidget_SAT_Room {
    label: "How Do Room Features Impact Lodging Satisfaction at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 2

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 85
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how room features, experiences and characteristics influence their overall lodging satisfaction. This shows us where to target improvement in our lodging processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT_EXPERIENCES.lodging
    independentVariables: surveyDataset:DRILL_ROOM.ac, surveyDataset:DRILL_ROOM.bathamenities, surveyDataset:DRILL_ROOM.bathclean, surveyDataset:DRILL_ROOM.bathfeatures, surveyDataset:DRILL_ROOM.bed, surveyDataset:DRILL_ROOM.cleanliness, surveyDataset:DRILL_ROOM.furnishings, surveyDataset:DRILL_ROOM.quiet, surveyDataset:DRILL_ROOM.smell, surveyDataset:DRILL_ROOM.wifi
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Room
  // widget keyDrivers #keyDriversWidget_SAT_Restaurants_Overall {
  //   label: "What Drives Restaurant Satisfaction Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 3 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }

  //   select #catfilter {
  //     label: "Filter by Meal Rated"
  //     mode: multi

  //     options: @categorySet_meal_rated.items
  //   }
  //   filter expression {
  //     value: selected(:MEAL_RATED, @catfilter.selected)
  //   }

    // algorithm: regression
    //// algorithm: correlation
  //   satisfactionLimit: 80
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
  //   importanceLimit: 0.15
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.restaurants
  //   independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Restaurants_Overall

  widget keyDrivers #keyDriversWidget_SAT_Restaurants {
    label: "What Drives Restaurant Satisfaction at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 3

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    select #catfilter {
      label: "Filter by Meal Rated"
      mode: multi

      options: @categorySet_meal_rated.items
    }
    filter expression {
      value: selected(:MEAL_RATED, @catfilter.selected)
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 80
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation

      size: large
    }
    description: "This analysis looks for patterns in the data to determine how different restaurant features influence their overall restaurant satisfaction. This shows us where to target improvement in our restaurant processes and experiences."
    importanceLimit: 0.15
    dependentVariable: surveyDataset:SAT_EXPERIENCES.restaurants
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Restaurants
  // widget keyDrivers #keyDriversWidget_SAT_Bars_Overall {
  //   label: "What Drives Bar Satisfaction Overall?"
  //   hide: @lodging_addl_keydrivers_selector.selected != 4 AND @Lodging_Locations_Selector.selected != "Lodging"

  //   // filter expression {
  //   //   value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

  //   // }

  //   scope reportingHierarchy {
  //     reportingHierarchy: SitesHierarchy
  //     nodes: AllData
  //   }
  //   minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    // algorithm: regression
    //// algorithm: correlation
  //   satisfactionLimit: 86
  //   showModelDetails: true
  //   quadrantTitles: @reportConfig.kda_quadrantTitles
  //   size: large
  //   infobox #infobox {
  //     label: @reportConfig.kda_infobox_label_correlation
  //     info: @reportConfig.kda_infobox_info_correlation
  //     size: large
  //   }
  //   description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the bar influence their overall bar satisfaction. This shows us where to target improvement in our bar processes and experiences."
  //   importanceLimit: 0.10
  //   dependentVariable: surveyDataset:SAT_EXPERIENCES.bars
  //   independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
  //   warningText: @reportConfig.kda_warningText
  // } // end widget keyDriversWidget_SAT_Bars_Overall

  widget keyDrivers #keyDriversWidget_SAT_Bars {
    label: "What Drives Bar Satisfaction at " + @Lodging_Locations_Selector.selectedLabel + "?"
    hide: @lodging_addl_keydrivers_selector.selected != 4

    filter expression {
      value: selected(:LocationFinal, @Lodging_Locations_Selector.selected)

    }

    scope reportingHierarchy {
      reportingHierarchy: SitesHierarchy
      nodes: AllData
    }

    minimumSampleSize: @reportConfig.KDAMinimumSampleSize
    algorithm: regression
    // algorithm: correlation

    defaultView: chart
    satisfactionLimit: 86
    showModelDetails: true
    quadrantTitles: @reportConfig.kda_quadrantTitles
    size: large
    infobox #infobox {
      label: @reportConfig.kda_infobox_label_regression
      info: @reportConfig.kda_infobox_info_regression

      // label: @reportConfig.kda_infobox_label_correlation
      // info: @reportConfig.kda_infobox_info_correlation
      size: large
    }
    description: "This analysis looks for patterns in the data to determine how aspects of a guest's experiences with the bar influence their overall bar satisfaction. This shows us where to target improvement in our bar processes and experiences."
    importanceLimit: 0.10
    dependentVariable: surveyDataset:SAT_EXPERIENCES.bars
    independentVariables: surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.quality
    warningText: @reportConfig.kda_warningText
  } // end widget keyDriversWidget_SAT_Bars
  widget headline #headlineWidget_17 {

    label: ""
    size: large

    tile markdown #markdownTile_2 {
      value: "## **Guest Comments**

### Comments provided by our guests represent the true voice of the customer - reviewing these comments can provide ideas for improvement and add clarity and context to the quantitative metrics shown in this report.

### Please note that you can select which comment to review (from the dropdown box); you can also sort  and filter the data that appears in each column."
    }

  } // end widget
  widget table #tableWidget {
    label: "Visitor Comments"
    size: "large"
    table: surveyDataset:

    showHeader: true
    sortOrder: descending
    sortColumn: comments

    headerNumberOfLines: 3
    stretchColumns: true

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response
    description: "This report shows specific comments guests made in the course of their feedback. To see more about a particular guest, please click the comment to show their full survey response."


    select #OpenEnd_selector {
      label: "Select Question"
      options: item {
        label: "Visit Comments"
        value:  {
          selectQuestion: surveyDataset:VISIT_COMMENTS
          selectFilter: surveyDataset:VISIT_COMMENTS != ""
        }

      },
      	    item {
        label: "Lodging Comments"
        value:  {
          selectQuestion: surveyDataset:LODGING_COMMENTS
          selectFilter: surveyDataset:LODGING_COMMENTS != ""
        }

      },
	    item {
        label: "Restaurant Comments"
        value:  {
          selectQuestion: surveyDataset:RESTAURANT_COMMENTS
          selectFilter: surveyDataset:RESTAURANT_COMMENTS != ""
        }

      },
      	    item {
        label: "Experiences Comments"
        value:  {
          selectQuestion: surveyDataset:EXPERIENCES_COMMENTS
          selectFilter: surveyDataset:EXPERIENCES_COMMENTS != ""
        }

      },
      item {
        label: "Problem Details"
        value:  {
          selectQuestion: surveyDataset:PROBLEM_DETAIL
          selectFilter: surveyDataset:PROBLEM_DETAIL != ""
        }

      },
      item {
        label: "Team Recognition"
        value:  {
          selectQuestion: surveyDataset:RECOG_DETAIL
          selectFilter: surveyDataset:RECOG_DETAIL != ""
        }

      }    

    } // end OpenEnd_selector
    filter expression {
      value: @OpenEnd_selector.selected.selectFilter
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }


    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }


    column response #comments {
      //sortBy: comment
      header: "Location: " + surveyDataset:LocationName
      footer: @reportConfig.intvdate
     // width: 300px
      enableColumnFilter: true
      comment: @OpenEnd_selector.selected.selectQuestion

    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Rec"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    column metric #copy_of_metricColumn {
      label: "OSAT"
      value: score(@reportConfig.osat_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

    column metric #copy_of_metricColumn2 {
      label: "Restaurants Sat"
      value: score(:DRILL_RESTAURANT.restaurant)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

  } // end widget

  widget headline #headlineWidget_15 {

    label: ""
    size: large
    hide: true
    tile markdown #markdownTile_2 {
      value: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    }

  }
  widget chart #chartWidget_NPS_Trends_Lines {
    label: "NPS® Trends"
    hide: true
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
    // ignoreFilters: reportingPeriod

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series1 {
      chart line {
        showDotValue: true

      }

      value: nps(@reportConfig.nps_qid) * 100
      format: noDecimalNumber
      label: "NPS®"

    }

    series #series2 {
      chart line {
        showDotValue: false

      }

      percentOver: series
      value: count(@reportConfig.nps_qid)
      format: oneDecimalPercent

      isSecondary: true
      breakdownBy cut {
        value: :NPSVal

      }
    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: noDecimalNumber
      label: "NPS®"
    }
    axis secondary #secondaryAxis {
      hide: false
      label: "% Response"
      format: noDecimalPercent
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      bottom: 75
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
  } // end widget
  widget chart #chartWidget_OSAT_Trends_Lines {
    label: "Overall Satisfaction (Top Box) Trend"
    // label: @kpiselect.selected.kpiLabel + " Trends"   
    palette: nps_and_cats_palette
    hide: true
    // ignoreFilters: reportingPeriod
    // hide: false

    // select #Timeframe_Selector {
    //   label: "Select Timeframe"

    //   options: @valueSet_date_ranges_1.items

    // } // end selector
    series #series1 {
      chart line {
        showDotValue: true

      }

      value: top1percent(@reportConfig.osat_qid)
      format: oneDecimalPercent
      label: "Overall Satisfaction"

    }

    category date #dateCategory {
      value: @reportConfig.intvdate
      breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
      label: "Interview date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      format: noDecimalPercent

    }
    axis primary #primaryAxis {
         //  format: metricsItemMetricDefaultFormatter
      format: oneDecimalPercent
      label: "Top Box % (5's)"
    }
    axis secondary #secondaryAxis {
      hide: true
      label: "% Response"
      format: noDecimalPercent
    }
    size: halfwidth

    legend: bottomCenter
    chartMargin {
      top: 20
      right: 20
      bottom: 75
    }

    base #base {
      value: count(@reportConfig.nps_qid)
      format: baseNumberFormatter
    }
    removeEmptyCategories: true
    removeEmptySeries: true
  } // end widget
  widget markdown #markdownWidget_PerformanceTrends {
    markdown: "# **Performance Trends**
### These tables provide a breakdown of how we perform on various key aspects of parks and resorts. In addition to Top Box scores (that is, the percentage of guests giving us the highest possible score), you can also see the monthly trend on each item."
    size: large
  }
  widget dataGrid #dataGridWidget_10 {
    label: "Satisfaction Drivers"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_DRIVERS$field
      total: none

    }
    column #column_current_counts {
      value: count(:SAT_DRIVERS$value)
      label: "Number of Responses"
      cell {
        value: count(:SAT_DRIVERS$value)
        format: noDecimalNumber
        //navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent
        //navigateTo: page_GamingResponses

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_DRIVERS$value)
        format: noDecimalPercent

        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }


  } //end widget
  widget dataGrid #dataGridWidget_ExperiencesSat {
    label: "Satisfaction with Experiences"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_EXPERIENCES$field
      total: none

    }
    column #column_current_counts {

      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:SAT_EXPERIENCES$value)

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell #undefined {
        format: noDecimalPercent
        value: top1percent(:SAT_EXPERIENCES$value)
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_EXPERIENCES$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_ResortExperiencesSat {
    label: "Satisfaction with Resort Experiences (Lizard)"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :SAT_RESORT_EXPERIENCES$field
      total: none

    }
    column #column_current_counts {

      label: "Number of Responses"
      cell #undefined {
        format: noDecimalNumber
        value: count(:SAT_RESORT_EXPERIENCES$value)

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell #undefined {
        format: noDecimalPercent
        value: top1percent(:SAT_RESORT_EXPERIENCES$value)
      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:SAT_RESORT_EXPERIENCES$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA

        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_LodgingSat {
    label: "Lodging Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_LODGING$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_LODGING$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_LODGING$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_LODGING$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RoomSat {
    label: "Room Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_ROOM$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_ROOM$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_ROOM$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_ROOM$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        //format: month
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
  widget dataGrid #dataGridWidget_RestaurantSat {
    label: "Restaurant Satisfaction"
    size: halfwidth
    removeEmptyColumns: true
    removeEmptyRows: true

    select #catfilter {
      label: "Filter by Meal Rated"
      mode: multi

      options: @categorySet_meal_rated.items
    }
    filter expression {
      value: selected(:MEAL_RATED, @catfilter.selected)
    }

    sort rows {
      sortBy: "/Satisfaction"
      sortOrder: descending
    }

    row cut {
      value: :DRILL_RESTAURANT$field
      total: none

    }
    column #column_current_counts {
      value: count(:DRILL_RESTAURANT$value)
      label: "Number of Responses"
      cell {
        value: count(:DRILL_RESTAURANT$value)
        format: noDecimalNumber

      }
    }

    column #column_Satisfaction {
      total: none
      label: "% Satisfied (Top Box)"
      cell {
        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent

      }
    }

    column #column_Satisfaction_Trends {
      label: "Satisfaction Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel

      cell microchart {

        value: top1percent(:DRILL_RESTAURANT$value)
        format: noDecimalPercent
        useOnlyExistingColumns: true
        breakdownBy date {
          value: @reportConfig.intvdate
          breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
        //format: month

        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } //end widget
//   widget headline #headlineWidget_LocationKPISummaries {

//     label: ""
//     size: large

//     tile markdown #markdownTile_2 {
//       value: "# **Location-Based KPI Summaries**
// ### This section looks at how specific locations track on our KPI's (and the trends)."
//     }

//   }
//   widget dataGrid #dataGridWidget_LocationPerfTrends {
//     label: "Location Performance Trends"
//     size: large
//     ignoreFilters: f_Location
//     removeEmptyRows: true

//     scope reportingHierarchy {
//       reportingHierarchy: SitesHierarchy
//       nodes: AllData
//     }

//     row comparison #comparisonRow {
//       reportingHierarchy: SitesHierarchySimplified
//       showTotal: false
//     }

//     column #column_Arrival {
//       label: "Arrival (Top Box)"
//       cell #cell {
//         value: top1percent(:DRILL_LODGING.arrival)
//         //target: @reportConfig.osat_target
//         format: oneDecimalPercent
//         extraValue: count(:DRILL_LODGING.arrival)
//         extraValueFormat: noDecimalNumber

//         navigateTo: page_LodgingResponses
//         navigateFilter: _isnotnull(:DRILL_LODGING.arrival)
//       }

//     }

//     column #column_Arrival_Trends {
//       label: "Arrival Sat Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
//       cell microchart #cell {
//         value: top1percent(:DRILL_LODGING.arrival)
//         format: oneDecimalPercent
//         useOnlyExistingColumns: true

//         microchart line #barMicrochart {
//           showDots: true
//           showTooltip: true
//           color: #1D78BA
//         }
//         breakdownBy date #dateBreakdownby {
//           value: @reportConfig.intvdate
//           breakdownBy: @Lodging_Timeframe_Selector.selected.selectBreakdownBy
//         //format: month

//         }
//       }

//     }

//     column #column_CleanRoom {
//       label: "Clean Room (Top Box)"
//       cell #cell {
//         value: top1percent(:DRILL_ROOM.cleanliness)
//         //target: @reportConfig.osat_target
//         format: oneDecimalPercent
//         extraValue: count(:DRILL_ROOM.cleanliness)
//         extraValueFormat: noDecimalNumber

//         navigateTo: page_LodgingResponses
//         navigateFilter: _isnotnull(:DRILL_ROOM.cleanliness)
//       }

//     }

//     column #column_CleanRoom_Trends {
//       label: "Clean Room Sat Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
//       cell microchart #cell {
//         value: top1percent(:DRILL_ROOM.cleanliness)
//         format: oneDecimalPercent
//         useOnlyExistingColumns: true

//         microchart line #barMicrochart {
//           showDots: true
//           showTooltip: true
//           color: #1D78BA
//         }
//         breakdownBy date #dateBreakdownby {
//           value: @reportConfig.intvdate
//           breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
//         //format: month

//         }
//       }

//     }

//     column #column_CleanBathroom {
//       label: "Clean Bathroom (Top Box)"
//       cell #cell {
//         value: top1percent(:DRILL_ROOM.bathclean)
//         //target: @reportConfig.osat_target
//         format: oneDecimalPercent
//         extraValue: count(:DRILL_ROOM.bathclean)
//         extraValueFormat: noDecimalNumber

//         navigateTo: page_LodgingResponses
//         navigateFilter: _isnotnull(:DRILL_ROOM.bathclean)
//       }

//     }

//     column #column_CleanBathroom_Trends {
//       label: "Clean Bathroom Sat Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
//       cell microchart #cell {
//         value: top1percent(:DRILL_ROOM.bathclean)
//         format: oneDecimalPercent
//         useOnlyExistingColumns: true

//         microchart line #barMicrochart {
//           showDots: true
//           showTooltip: true
//           color: #1D78BA
//         }
//         breakdownBy date #dateBreakdownby {
//           value: @reportConfig.intvdate
//           breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
//         //format: month

//         }
//       }

//     }

//     column #column_Restaurants {
//       label: "Restaurants Sat (Top Box)"
//       cell #cell {
//         value: top1percent(:SAT_EXPERIENCES.restaurants)
//         //target: @reportConfig.osat_target
//         format: oneDecimalPercent
//         extraValue: count(:SAT_EXPERIENCES.restaurants)
//         extraValueFormat: noDecimalNumber

//         navigateTo: page_LodgingResponses
//         navigateFilter: _isnotnull(:SAT_EXPERIENCES.restaurants)
//       }

//     }
//     column #column_Restaurants_Trends {
//       label: "Restaurants Sat Trends" + " - " + @Australia_Timeframe_Selector.selectedLabel
//       cell microchart #cell {
//         value: top1percent(:SAT_EXPERIENCES.restaurants)
//         format: oneDecimalPercent
//         useOnlyExistingColumns: true

//         microchart line #barMicrochart {
//           showDots: true
//           showTooltip: true
//           color: #1D78BA
//         }
//         breakdownBy date #dateBreakdownby {
//           value: @reportConfig.intvdate
//           breakdownBy: @Australia_Timeframe_Selector.selected.selectBreakdownBy
//         //format: month

//         }
//       }

//     }

//     infobox #infobox {
//       label: "Sites KPIs info"
//       info: ""
//     }
//     showLegend: true
//     view comparativeStatistic #comparativeStatisticView {
//       valueColorFormatter: copy_of_sentimentindicatortext
//       backgroundColorFormatter: gridDefaultBackgroundColorFormatter
//     }
//   } // end widget
  //hide: false
  modal: false
} // end page
page #page_CasesOverview {
  label: "Action Management"

  access rules {
    rule claim {
      name: "UserLevel"
      value: "Power User", "Field"
    }
  }

  layoutArea toolbar {
  //useDynamicFilters: true

  } // end page layoutArea
  widget headline #totalOpenCases {
    label: "All ʺOpenʺ cases"


    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOpen()
      label: "Cases - Open"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: openCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOpenʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #copy_of_totalOpenCases {
    label: "All ʺIn Progressʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesInProg()
      label: "Cases - In Progress"
    }

    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: inprogressCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺIn-Progressʺ and need attention."
      fontSize: 20
    }

  } // end widget
  widget headline #totalInProgressCases {
    label: "All ʺOverdueʺ cases"

    filter expression #expressionFilter {
      value: amTable:filterMeasure_AMCasesOverdue()
      label: "Cases - Overdue"
    }
    tile value #valueTile {
      value: count(amTable:CaseId)
      fontSize: 129
      valueColorFormatter: overdueCasesColorFormatter_1
    }

    tile text #textTile {
      value: "These alerts are ʺOverdueʺ and need attention."
      fontSize: 20
    }
  } // end widget
  widget chart #daystoClose {

    label: "Average Days To Close"
    size: halfwidth
    gridLines: horizontal
    removeEmptyCategories: true

    filter expression {
      value: amTable:SystemStatus = "closed"
    }

    chartMargin {
      right: 60
      bottom: 50
    }
    chart area {
      lineType: monotone

    }

    series {
      label: "Average Days to Close"
      value: median(amTable:daysToClose)
    }

    category cut {
      value: amTable:Workflow
    }

    axis primary #primaryAxis {
      axisLine: true
      tickLine: true
    }
    axis category #categoryAxis {
      axis secondary #secondaryAxis {
        hide: true
      }
      orientation: "-45"
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    removeEmptySeries: true
  } //end widget
  widget chart #topCXissues {
    label: "Top Case Types"
    gridLines: horizontal
    removeEmptySeries: true
    removeEmptyCategories: true
    size: halfwidth

    chartMargin {
      right: 60
      bottom: 50
    }

    series #series {
      chart bar #barChart {
        maxBarSize: 50
      }
      value: count(amTable:Trigger)
    }

    axis primary #primaryAxis {
      axisLine: true
      tickLine: true
      minValue: 0
      maxValue: -1
    }
    category cut #cutCategory {
      value: amTable:Trigger
    }

    axis secondary #secondaryAxis {
      hide: true
    }
    axis category #categoryAxis {
      orientation: "-45"
    }
  } //end widget
  widget table #tableWidget {
    label: "Cases"
    size: "large"
    table: amTable:
    sortColumn: DateCreated
    sortOrder: descending
    paginationType: paging
    rowsPerPage: 100,150,250,500
    navigateTo: page_CaseDetails


    view metric #metricView {
      backgroundColorFormatter: TableBackgroundColorFormatter
      valueColorFormatter: dropOffDefaultFormatter
    }

    column date #DateCreated {
      label: "Date Created"
      value: amTable:DateCreated
      enableColumnFilter: true
    }

    column value #location {
      label: "Location"
      value: surveyDataset:LocationName
      sortable: true
      enableColumnFilter: true
    }

    column value #CaseId {
      label: "CaseId"
      value: amTable:CaseId
      enableColumnFilter: true
    }

    column value #caseStatus {
      label: "Case Status"
      value: amTable:lk_3827
      enableColumnFilter: true
    }

    column value #valueColumn_4 {
      label: "Case Name"
      value: amTable:CaseName
      enableColumnFilter: true
    }
    column value #guestname {
      label: "Guest Name"
      value: surveyDataset:guest_name
      sortable: true
      enableColumnFilter: true
    }
    column value #rank_description {
      label: "Lucky North tier designation"
      value: surveyDataset:rank_description
      sortable: true
      enableColumnFilter: true
    }

    column value #team_member {
      label: "Team Member"
      value: surveyDataset:TEAM_MEMBER
      sortable: true
      enableColumnFilter: true
    }
    column value #recog_comments {
      label: "Recognition Comments"
      value: surveyDataset:RECOG_DETAIL
      sortable: true
      enableColumnFilter: true
    }

    column value #problem_comments {
      label: "Problem Comments"
      value: surveyDataset:PROBLEM_DETAIL
      sortable: true
      enableColumnFilter: true
    }

    column value #visit_comments {
      label: "Visit Comments"
      value: surveyDataset:VISIT_COMMENTS
      sortable: true
      enableColumnFilter: true
    }

  } //end widget
} // end page
page #page_CaseDetails {
  label: "Case Details"
  layoutArea toolbar {
    hide: true
  }
  hide: true
  widget caseDetailsSummary {
    size: large
  }
  widget caseResponse {
    size: halfwidth
    showSegmentedBars: true
    hideUnansweredDefault: true
  }
  widget caseManagement {
    size: halfwidth
  }
  widget caseLog {
    size: large
  }
} // end page
page #page_NPSResponses {
  label: "NPS Responses"
  modal: true
  widget table #tableWidget {
    label: "NPS Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start
    rowsPerPage: 100, 500, 1000

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: large
    }

    view metric #colorcoding_11pt {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    filter expression {
      value: surveyDataset:filterMeasure_NPSanswered()
      label: "NPS has a value"
    }

    column value #SurveyName {
      label: "Survey"
      value: surveyDataset:survey_pid
      enableColumnFilter: true
      align: center
      width: 100px

    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
      align: center
      width: 100px
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
      align: center
      width: 100px
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
      align: center
      width: 50px
    }


    column value #LocationName {
      label: "Location"
      //value: demote(SitesHierarchy:language_text, surveyDataset:)
      value: surveyDataset:LocationName
      enableColumnFilter: true
      align: center
      width: 200px
    }

    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 100px
      align: center
      enableColumnFilter: true
    }

    column metric #metricColumn {
      label: "Likely to Rec"
      value: @reportConfig.nps_qid
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_11pt

    }
    column metric #copy_of_metricColumn {
      label: "OSAT"
      value: score(@reportConfig.osat_qid)
      enableColumnFilter: true
      width: 100px
      align: center
      view: colorcoding_5pt

    }

    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
          //  align: center
      width: 200px
    }

    navigateTo: page_Indiv_Survey_Response
  } // end widget
} // end page
page #page_Responses_modal {
  label: "Responses"
  //modal: true

  widget table #ResponsesTable_Modal {
    label: "Responses"
    table: :
    size: halfwidth

    sortColumn: ResponseDate
    sortOrder: descending
    paginationType: paging
    rowsPerPage: 50, 100, 250

    filter expression {
      value: _isnotnull(@reportConfig.nps_qid)
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2 //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: small
    }

    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: small
    }

    column date #ResponseDate {
      label: "Response Date"
      value: :interview_start
      format: dateDefaultFormatter
      //format: dateFormatDay

      enableColumnFilter: true
      align: center
      width: 50px
    }

    column value #SurveyName {
      label: "Survey"
      value: surveyDataset:survey_pid
      enableColumnFilter: true
      align: center
      width: 50px

    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset:LocationName
      enableColumnFilter: true
      align: center
      width: 50px

    }


    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 50px
      align: center
      enableColumnFilter: true
    }

    column metric #nps {
      label: "NPS"
      value: @reportConfig.nps_qid
      align: center
      //format: colorFormatter
      view: colorcoding
      width: 50px
      enableColumnFilter: true
    }
    column value #comments {
      label: "Visit Comments"
      value: surveyDataset:VISIT_COMMENTS
      width: 100px
      enableColumnFilter: true

    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
    }

    navigateTo: page_Indiv_Survey_Response
  } // end widget
  config layout #layoutConfig {
    horizontalAlignmentMode: "fullWidth"
  }

  hide: false
  modal: true
  modalSize: large
} // end page
page #page_Problem_Responses_modal {
  label: "Problem Responses"
  //modal: true

  widget table #ResponsesTable_Modal {
    label: "Responses"
    table: :
    size: halfwidth

    sortColumn: ResponseDate
    sortOrder: descending
    paginationType: paging
    rowsPerPage: 50, 100, 250

    filter expression {
      value: _isnotnull(@reportConfig.nps_qid)
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2 //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: small
    }

    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: small
    }

    column date #ResponseDate {
      label: "Response Date"
      value: :interview_start
      format: dateDefaultFormatter
      //format: dateFormatDay

      enableColumnFilter: true
      align: center
      width: 50px
    }

    column value #SurveyName {
      label: "Survey"
      value: surveyDataset:survey_name
      enableColumnFilter: true
      align: center
      width: 50px

    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset:LocationName
      enableColumnFilter: true
      align: center
      width: 50px

    }


    column metric #metricColumn_1 {
      label: "NPS Segment"
      value: score(surveyDataset:NPSVal)
      format: npssegmentindicatortextValue2
      target: 9
      view: viewnpssegment
      width: 50px
      align: center
      enableColumnFilter: true
    }

    column metric #nps {
      label: "NPS"
      value: @reportConfig.nps_qid
      align: center
      //format: colorFormatter
      view: colorcoding
      width: 30px
      enableColumnFilter: true
    }


    column value #valueColumn_4 {
      label: "Problem"
      value: :PROBLEM
      width: 50px
      enableColumnFilter: true
    }
    column value #valueColumn_5 {
      label: "Problem Details"
      value: :PROBLEM_DETAIL
      width: 100px
      enableColumnFilter: true
    }
    column value #valueColumn_6 {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      width: 30px
      enableColumnFilter: true
    }
    column value #valueColumn_7 {
      label: "Problem Reported"
      value: :PROB_REPORTED
      width: 30px
      enableColumnFilter: true
    }
    navigateTo: page_Indiv_Survey_Response
  } // end widget
  config layout #layoutConfig {
    horizontalAlignmentMode: "fullWidth"
  }

  hide: false
  modal: true
  modalSize: large
} // end page
page #page_ProblemDrilldown {
  label: "Problem Drill-Down"
  widget table #tableWidget {
    label: "Guests Requesting Contact"
    size: "large"
    table: :
    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_ContactRequested()
      label: "Contact Req = Yes"
    }

    column value #valueColumn_7 {
      label: "Location"
      value: :LocationName
      enableColumnFilter: true
    }
    column value #valueColumn {
      label: "Guest Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "Guest Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #valueColumn_3 {
      label: "Guest Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #valueColumn_4 {
      label: "Contact Preference"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #valueColumn_5 {
      label: "Guest Notes on Problem"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #valueColumn_6 {
      label: "Sat with Problem Resolution"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    navigateTo: page_Indiv_Survey_Response
  } //end widget
  widget chart #chartWidget_3 {
    label: "Problem During Visit?"
    series #series {
      value: count(:PROBLEM)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
      //navigateTo: page_ProblemDrilldown
      //navigateFilter: surveyDataset:filterMeasure_DNListensSurvey()
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: small
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomCenter"


    category cut #cutCategory {
      value: :PROBLEM

    }
    palette: redtogreen2ptscale
  } //end widget
  widget chart #copy_of_chartWidget_4 {
    label: "Problem Reported?"
    series #series {
      value: count(:respid)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: large
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomLeft"
    category cut #cutCategory {
      value: :PROB_REPORTED
    }
    palette: redtogreen2ptscale
  }
  widget kpi #kpiWidget {
    label: "Satisfaction with Problem Resolution"
    size: small
    tile kpi #kpiTile {
      value: top1percent(:RESOLUTION_SAT)
      //  value: 35
      label: "Resolution SAT (5's)"

      format: percentDefaultFormatter
      min: 0
      max: 100

      targetFormat: noDecimalNumber
      showRange: true
      belowTargetLabel: @reportConfig.belowTargetLabel
      aboveTargetLabel: @reportConfig.aboveTargetLabel
      atTargetLabel: @reportConfig.atTargetLabel
    }

    tile value #valueTile {
      value: count(:RESOLUTION_SAT)
      label: "Responses"
      format: noDecimalNumber
    }
    //description: "This shows our Overall Satisfaction KPI, which is based on the extent to which guests are ʺVery Satisfiedʺ with their entire experience. To see more information on Overall Satisfaction, please click the ʺiʺ icon above."
    tile value #valueTile_2 {
      value: average(numeric(:RESOLUTION_SAT))
      label: "Average Satisfaction Score"
      min: 1
      max: 5
    }
    tile value #valueTile_3 {
      value: bottom2percent(:RESOLUTION_SAT)
      label: "% Dissatisfied"
      min: 0
      max: 100
      format: percentDefaultFormatter
    }
  } //end widget
  widget chart #copy_of_copy_of_chartWidget_4 {
    label: "Would You Like to be Contacted?"
    series #series {
      value: count(:respid)
      format: percentDefaultFormatter
      chart pie #pieChart {
        showBase: true
      }
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: large
    chart pie #pieChart {
      legendType: square
    }
    legend: "bottomLeft"
    category cut #cutCategory {
      value: :CONTACT
    }
    palette: redtogreen2ptscale
  } //end widget
  hide: false
  modal: true
  modalSize: "large"
} // end page
page #page_TeamRecog {
  label: "Team Member Recognition"
  widget table #tableWidget {
    label: "Recognition from Guests"
    size: "large"
    table: :

    column value #valueColumn_7 {
      label: "Location"
      value: :LocationName
      enableColumnFilter: true
    }
    column value #valueColumn {
      label: "Team Member Name"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #valueColumn_4 {
      label: "Guest Recognition Notes"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }
    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_TeamRecog()
      label: "Recog = Yes"
    }
    navigateTo: page_Indiv_Survey_Response
  }
  hide: false
  modal: true
  modalSize: "large"
} // end page
page #page_Indiv_Survey_Response {
  label: "Individual Survey Response"
  widget contactSurveyResponse #contactSurveyResponseWidget {
    label: "Individual Survey Response"

    config individualResponse #individualResponseConfig {
      summary #summary {
        variables: surveyDataset:survey_name, surveyDataset:survey_rid, surveyDataset:LocationName
      }

      tab #tab_survey_data {
        tile list #listTile {
          variables: surveyDataset:interview_start, surveyDataset:status, surveyDataset:SurveyType, surveyDataset:LocationName, surveyDataset:VISIT_DATE, surveyDataset:TIME_OF_VISIT, surveyDataset:STORE_INFO, surveyDataset:LocationWeb, surveyDataset:StateProvince, surveyDataset:NPS, surveyDataset:RETURN_VISIT, surveyDataset:SAT, surveyDataset:GAMING_EXPERIENCES, surveyDataset:GamingSurveyPath, surveyDataset:Value, surveyDataset:EXPERIENCES, surveyDataset:EXP_DRILLFLAG, surveyDataset:SAT_DRIVERS.staff, surveyDataset:SAT_DRIVERS.cleanliness, surveyDataset:SAT_DRIVERS.eodb, surveyDataset:SAT_DRIVERS.safety, surveyDataset:SAT_DRIVERS.quality, surveyDataset:SAT_DRIVERS.value, surveyDataset:SAT_DRIVERS.variety, surveyDataset:SAT_DRIVERS.speed, surveyDataset:EDUC_EXP.educational, surveyDataset:SAT_GAMING.gaming, surveyDataset:SAT_GAMING.playersclub, surveyDataset:SAT_GAMING.pokerroom, surveyDataset:SAT_GAMING.slots, surveyDataset:SAT_GAMING.tablegames, surveyDataset:SAT_GAMING.betting, surveyDataset:SAT_GAMING.drinks, surveyDataset:SAT_GAMING.restaurants, surveyDataset:SAT_GAMING.bars, surveyDataset:SAT_GAMING.buffet, surveyDataset:SAT_GAMING.lodging, surveyDataset:VISIT_COMMENTS, surveyDataset:TICKETS, surveyDataset:PURPOSE_VISIT, surveyDataset:ARRIVAL.1, surveyDataset:ARRIVAL.2, surveyDataset:ARRIVAL.3, surveyDataset:ARRIVAL.4, surveyDataset:ARRIVAL.5, surveyDataset:ARRIVAL.6, surveyDataset:SAT_EXPERIENCES.attractions, surveyDataset:SAT_EXPERIENCES.bus, surveyDataset:SAT_EXPERIENCES.restaurants, surveyDataset:SAT_EXPERIENCES.premiums, surveyDataset:SAT_EXPERIENCES.shops, surveyDataset:SAT_EXPERIENCES.rides, surveyDataset:SAT_EXPERIENCES.breakfast, surveyDataset:SAT_EXPERIENCES.bars, surveyDataset:SAT_EXPERIENCES.concierge, surveyDataset:SAT_EXPERIENCES.spa, surveyDataset:SAT_EXPERIENCES.otheramenities, surveyDataset:ATTRACTIONS_SEEN, surveyDataset:ATTRACT_INSERT, surveyDataset:DRILL_ATTRACTION.quality, surveyDataset:DRILL_ATTRACTION.cleanliness, surveyDataset:DRILL_ATTRACTION.staff, surveyDataset:DRILL_BUS.quality, surveyDataset:DRILL_BUS.staff, surveyDataset:DRILL_BUS.waitime, surveyDataset:DRILL_BUS.cleanarea, surveyDataset:DRILL_BUS.cleanbus, surveyDataset:DRILL_SLOTS.selection, surveyDataset:DRILL_SLOTS.avail, surveyDataset:DRILL_TABLEGAMES.selection, surveyDataset:DRILL_TABLEGAMES.betting, surveyDataset:DRILL_TABLEGAMES.avail, surveyDataset:DRILL_TABLEGAMES.staff, surveyDataset:DRILL_GAME_DRINK.value, surveyDataset:DRILL_GAME_DRINK.speed, surveyDataset:DRILL_GAME_DRINK.taste, surveyDataset:DRILL_LODGING.accuracy, surveyDataset:DRILL_LODGING.arrival, surveyDataset:DRILL_LODGING.cleanliness, surveyDataset:DRILL_LODGING.avail, surveyDataset:DRILL_LODGING.staff, surveyDataset:DRILL_LODGING.service, surveyDataset:DRILL_LODGING.departure, surveyDataset:DRILL_ROOM.cleanliness, surveyDataset:DRILL_ROOM.furnishings, surveyDataset:DRILL_ROOM.ac, surveyDataset:DRILL_ROOM.smell, surveyDataset:DRILL_ROOM.quiet, surveyDataset:DRILL_ROOM.bed, surveyDataset:DRILL_ROOM.wifi, surveyDataset:DRILL_ROOM.bathclean, surveyDataset:DRILL_ROOM.bathfeatures, surveyDataset:DRILL_ROOM.bathamenities, surveyDataset:LODGING_COMMENTS, surveyDataset:ROOM_COMMENTS, surveyDataset:RESTAURANT_INSERT_TEXT, surveyDataset:MEAL_RATED, surveyDataset:DRILL_RESTAURANT.quality, surveyDataset:DRILL_RESTAURANT.value, surveyDataset:DRILL_RESTAURANT.staff, surveyDataset:DRILL_RESTAURANT.kiosk, surveyDataset:DRILL_RESTAURANT.speed, surveyDataset:DRILL_RESTAURANT.variety, surveyDataset:DRILL_RESTAURANT.cleanliness, surveyDataset:DRILL_BUFFET.quality, surveyDataset:DRILL_BUFFET.value, surveyDataset:DRILL_BUFFET.variety, surveyDataset:DRILL_BUFFET.stock, surveyDataset:DRILL_BUFFET.taste, surveyDataset:DRILL_BUFFET.temperature, surveyDataset:DRILL_BUFFET.cleanliness, surveyDataset:DINING_COMMENT_INSERT, surveyDataset:RESTAURANT_COMMENTS, surveyDataset:PREMIUM_PURCHASED, surveyDataset:PREMIUM_INSERT, surveyDataset:DRILL_PREMIUM.quality, surveyDataset:DRILL_PREMIUM.value, surveyDataset:DRILL_PREMIUM.staff, surveyDataset:DRILL_PREMIUM.foodquality, surveyDataset:SHOPS_VISITED, surveyDataset:SHOPS_INSERT, surveyDataset:PURCHASE, surveyDataset:DRILL_SHOPS.shopsat, surveyDataset:DRILL_SHOPS.value, surveyDataset:DRILL_SHOPS.staff, surveyDataset:DRILL_SHOPS.speed, surveyDataset:DRILL_SHOPS.merch, surveyDataset:DRILL_SHOPS.variety, surveyDataset:BOOKING_METHOD, surveyDataset:DRILL_BOOKING.bookingsat, surveyDataset:DRILL_BOOKING.avail, surveyDataset:DRILL_BOOKING.info, surveyDataset:DRILL_BOOKING.communication, surveyDataset:BOOKING_COMMENTS, surveyDataset:DRILL_TOURS.avail, surveyDataset:DRILL_TOURS.staff, surveyDataset:DRILL_TOURS.knowledge, surveyDataset:DRILL_TOURS.equipment, surveyDataset:TOURS_COMMENTS, surveyDataset:TOURS_ELEMENTS.guidesat, surveyDataset:TOURS_ELEMENTS.knowledge, surveyDataset:TOURS_ELEMENTS.toursafety, surveyDataset:TOURS_ELEMENTS.sitesat, surveyDataset:TOURS_ELEMENTS.cleanbus, surveyDataset:TOURS_ELEMENTS.lunch, surveyDataset:ELEMENTS_COMMENT, surveyDataset:PROBLEM, surveyDataset:PROB_REPORTED, surveyDataset:RESOLUTION_SAT, surveyDataset:CONTACT, surveyDataset:CONTACT_PREF, surveyDataset:CONTACT_INFO.name, surveyDataset:CONTACT_INFO.phone, surveyDataset:CONTACT_INFO.email, surveyDataset:PROBLEM_DETAIL, surveyDataset:TEAM_REC, surveyDataset:TEAM_MEMBER, surveyDataset:RECOG_DETAIL, surveyDataset:REGION, surveyDataset:GENDER, surveyDataset:AGE, surveyDataset:INCOME, surveyDataset:UNDER_18_KIDS, surveyDataset:EDUCATION, surveyDataset:ETHNICITY, surveyDataset:COMPANIONS, surveyDataset:TOTAL_PARTY, surveyDataset:TIME_OF_GAMING_VISIT, surveyDataset:WIN_LOSE, surveyDataset:SPEC_EVENT, surveyDataset:COMPS, surveyDataset:REDEMPTION, surveyDataset:NO_VISITS, surveyDataset:AWARENESS, surveyDataset:KSC_COMPANIONS, surveyDataset:ACCOMMODATIONS, surveyDataset:LOCATION, surveyDataset:OTHER_ATTRACTIONS, surveyDataset:NO_VACATIONS, surveyDataset:LOI, surveyDataset:Southland_Gaming_Seg_assign, surveyDataset:Southland_Gaming_Seg_scores.1, surveyDataset:Southland_Gaming_Seg_scores.2, surveyDataset:Southland_Gaming_Seg_scores.3, surveyDataset:Southland_Gaming_Seg_scores.4, surveyDataset:Southland_Gaming_Seg_scores.5, surveyDataset:GAMING_SEGMENTATION.funexperience, surveyDataset:GAMING_SEGMENTATION.winagain, surveyDataset:GAMING_SEGMENTATION.relax, surveyDataset:GAMING_SEGMENTATION.entertain, surveyDataset:GAMING_SEGMENTATION.lifechanging, surveyDataset:GAMING_SEGMENTATION.overnightstay, surveyDataset:GAMING_SEGMENTATION.skills, surveyDataset:GAMING_SEGMENTATION.funalone, surveyDataset:GAMING_SEGMENTATION.tobesurprised, surveyDataset:GAMING_SEGMENTATION.treatmyself
        }
        label: "Survey Results"
      }


      tab #tab_BG_info {
        tile list #listTile {
          variables: surveyDataset:LocationName, surveyDataset:email, surveyDataset:customer_id, surveyDataset:player_id, surveyDataset:guest_name, surveyDataset:guest_gender, surveyDataset:customer_state, surveyDataset:Postal, surveyDataset:customer_country, surveyDataset:customer_city, surveyDataset:date_of_birth, surveyDataset:guest_age, surveyDataset:TransactionID, surveyDataset:transaction_time_stamp, surveyDataset:YieldDateTime, surveyDataset:CountryName, surveyDataset:CompanyID, surveyDataset:NodeNo, surveyDataset:SellingPrice, surveyDataset:UseNo, surveyDataset:visits, surveyDataset:minutes_played, surveyDataset:avgADT, surveyDataset:game_pref, surveyDataset:rank_description, surveyDataset:last_play_date, surveyDataset:date_enrolled, surveyDataset:total_guest_count, surveyDataset:children_count, surveyDataset:adult_count, surveyDataset:reservation_revenue, surveyDataset:market_segment_code, surveyDataset:reservation_status, surveyDataset:room_description, surveyDataset:room_category, surveyDataset:rate_description, surveyDataset:departure_date, surveyDataset:arrival_date, surveyDataset:confirm_number
        }
        label: "Background Info"
      }

    }
    size: halfwidth
    table: :
    showUnanswered: false
    view bar #surveyResponseItemBarDefaultView {
      chartColorFormat: scoreNPS_blue
    }
  } //end widget
  hide: false
  modal: true
} // end page
page #page_Indiv_Survey_Response_TA {
  label: "Individual Survey Response-TA"
  widget contactSurveyResponse #contactSurveyResponseWidget {
    label: "Individual Survey Response"

    config individualResponse #individualResponseConfig {
      summary #summary {
        variables: surveyDataset_TA:survey_name, surveyDataset_TA:LocationName, surveyDataset_TA:rank_description, surveyDataset_TA:interview_start, surveyDataset_TA:status
      }

      tab #tab_survey_data {
        tile list #listTile {
          variables: surveyDataset_TA:survey_rid, surveyDataset_TA:VISIT_DATE, surveyDataset_TA:STORE_INFO, surveyDataset_TA:NPS, surveyDataset_TA:SAT, surveyDataset_TA:Value, surveyDataset_TA:VISIT_COMMENTS_DNLISTENS, surveyDataset_TA:VISIT_COMMENTS_KSCVC, surveyDataset_TA:VISIT_COMMENTS_LODGING, surveyDataset_TA:VISIT_COMMENTS_GAMING, surveyDataset_TA:VISIT_COMMENTS_TOURS, surveyDataset_TA:VISIT_COMMENTS_LIZARD, surveyDataset_TA:LODGING_COMMENTS_LODGING, surveyDataset_TA:LODGING_COMMENTS_GAMING, surveyDataset_TA:LODGING_COMMENTS_LIZARD, surveyDataset_TA:ROOM_COMMENTS_LODGING, surveyDataset_TA:RESTAURANT_COMMENTS_KSCVC, surveyDataset_TA:RESTAURANT_COMMENTS_LODGING, surveyDataset_TA:RESTAURANT_COMMENTS_GAMING, surveyDataset_TA:RESTAURANT_COMMENTS_LIZARD, surveyDataset_TA:BOOKING_COMMENTS_TOURS, surveyDataset_TA:TOURS_COMMENTS, surveyDataset_TA:ELEMENTS_COMMENT_TOURS, surveyDataset_TA:EXPERIENCES_COMMENTS_LIZARD, surveyDataset_TA:PROBLEM,  surveyDataset_TA:PROB_REPORTED,  surveyDataset_TA:RESOLUTION_SAT, surveyDataset_TA:PROBLEM_DETAIL_DNLISTENS, surveyDataset_TA:PROBLEM_DETAIL_KSCVC, surveyDataset_TA:PROBLEM_DETAIL_LODGING, surveyDataset_TA:PROBLEM_DETAIL_GAMING, surveyDataset_TA:PROBLEM_DETAIL_LIZARD, surveyDataset_TA:TEAM_REC, surveyDataset_TA:TEAM_MEMBER, surveyDataset_TA:RECOG_DETAIL_DNLISTENS, surveyDataset_TA:RECOG_DETAIL_KSCVC, surveyDataset_TA:RECOG_DETAIL_LODGING, surveyDataset_TA:RECOG_DETAIL_GAMING, surveyDataset_TA:RECOG_DETAIL_LIZARD
        }
        label: "Survey Results"
      }

      tab #tab_demos_data {
        tile list #listTile {
          variables: surveyDataset_TA:REGION, surveyDataset_TA:REGION_ALPHA, surveyDataset_TA:GENDER, surveyDataset_TA:AGE, surveyDataset_TA:INCOME, surveyDataset_TA:UNDER_18_KIDS, surveyDataset_TA:EDUCATION, surveyDataset_TA:ETHNICITY, surveyDataset_TA:ETHNICITY_AUS
        }
        label: "Demographics"
      }


      tab #tab_BG_info {
        tile list #listTile {
          variables: surveyDataset_TA:LocationName, surveyDataset_TA:TransactionID, surveyDataset_TA:guest_name, surveyDataset_TA:rank_description
        }
        label: "Background Info"
      }

    }
    size: halfwidth
    table: surveyDataset_TA:
    showUnanswered: false
    view bar #surveyResponseItemBarDefaultView {
      chartColorFormat: scoreNPS_blue
    }
  } //end widget
  hide: false
  modal: true
} // end page
page #page_ResponseDetails {

  label: "Response Details"

  access rules {
    rule claim {
      name: "UserLevel"
      value: "Power User"
    }
  }

  widget table #tableWidget {
    label: "Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start
    rowsPerPage: 100, 500, 1000

    column value #SurveyName {
      label: "Survey Name"
      value: :survey_pid
      enableColumnFilter: true
    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
    }

    column value #SurveyType {
      label: "Survey Type (DN Listens)"
      value: :SurveyType
      enableColumnFilter: true
    }
    column value #LocationName {
      label: "Location Name"
      value: :LocationName
      enableColumnFilter: true
    }
    column date #VISIT_DATE {
      label: "Visit Date"
      value: :VISIT_DATE
      enableColumnFilter: true
    }
    column value #TIME_OF_VISIT {
      label: "Time of Visit"
      value: :TIME_OF_VISIT
      enableColumnFilter: true
    }
    column value #STORE_INFO {
      label: "Store Info"
      value: :STORE_INFO
      enableColumnFilter: true
    }
    // column value #valueColumn_8 {
    //   label: "LocationWeb"
    //   value: :LocationWeb
    //   enableColumnFilter: true
    // }
    column value #StateProvince {
      label: "State / Province"
      value: :StateProvince
      enableColumnFilter: true
    }
    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
    }

    column value #RETURN_VISIT {
      label: "Return Visit"
      value: :RETURN_VISIT
      enableColumnFilter: true
    }
    column value #SAT {
      label: "SAT"
      value: :SAT
      enableColumnFilter: true
    }
    column value #GAMING_EXPERIENCES {
      label: "GAMING_EXPERIENCES"
      value: :GAMING_EXPERIENCES
      enableColumnFilter: true
    }
    column value #GamingSurveyPath {
      label: "GamingSurveyPath"
      value: :GamingSurveyPath
      enableColumnFilter: true
    }
    column value #Value {
      label: "Value"
      value: :Value
      enableColumnFilter: true
    }
    column value #EXPERIENCES {
      label: "EXPERIENCES"
      value: :EXPERIENCES
      enableColumnFilter: true
    }
    column value #EXP_DRILLFLAG {
      label: "EXP_DRILLFLAG"
      value: :EXP_DRILLFLAG
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_cleanliness {
      label: "SAT_DRIVERS.cleanliness"
      value: :SAT_DRIVERS.cleanliness
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_eodb {
      label: "SAT_DRIVERS.eodb"
      value: :SAT_DRIVERS.eodb
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_quality {
      label: "Food quality"
      value: :SAT_DRIVERS.quality
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_safety {
      label: "SAT_DRIVERS.safety"
      value: :SAT_DRIVERS.safety
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_speed {
      label: "Speed of service"
      value: :SAT_DRIVERS.speed
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_staff {
      label: "Staff"
      value: :SAT_DRIVERS.staff
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_value {
      label: "Value"
      value: :SAT_DRIVERS.value
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_variety {
      label: "Variety of items"
      value: :SAT_DRIVERS.variety
      enableColumnFilter: true
    }
    column value #EDUC_EXP {
      label: "EDUC_EXP.educational"
      value: :EDUC_EXP.educational
      enableColumnFilter: true
    }
    column value #SAT_GAMING_bars {
      label: "SAT_GAMING.bars"
      value: :SAT_GAMING.bars
      enableColumnFilter: true
    }
    column value #SAT_GAMING_betting {
      label: "SAT_GAMING.betting"
      value: :SAT_GAMING.betting
      enableColumnFilter: true
    }
    column value #SAT_GAMING_buffet {
      label: "SAT_GAMING.buffet"
      value: :SAT_GAMING.buffet
      enableColumnFilter: true
    }
    column value #SAT_GAMING_drinks {
      label: "SAT_GAMING.drinks"
      value: :SAT_GAMING.drinks
      enableColumnFilter: true
    }
    column value #SAT_GAMING_gaming {
      label: "SAT_GAMING.gaming"
      value: :SAT_GAMING.gaming
      enableColumnFilter: true
    }
    column value #SAT_GAMING_lodging {
      label: "SAT_GAMING.lodging"
      value: :SAT_GAMING.lodging
      enableColumnFilter: true
    }
    column value #SAT_GAMING_playersclub {
      label: "SAT_GAMING.playersclub"
      value: :SAT_GAMING.playersclub
      enableColumnFilter: true
    }
    column value #SAT_GAMING_pokerroom {
      label: "SAT_GAMING.pokerroom"
      value: :SAT_GAMING.pokerroom
      enableColumnFilter: true
    }
    column value #SAT_GAMING_restaurants {
      label: "SAT_GAMING.restaurants"
      value: :SAT_GAMING.restaurants
      enableColumnFilter: true
    }
    column value #SAT_GAMING_slots {
      label: "SAT_GAMING.slots"
      value: :SAT_GAMING.slots
      enableColumnFilter: true
    }
    column value #SAT_GAMING_tablegames {
      label: "SAT_GAMING.tablegames"
      value: :SAT_GAMING.tablegames
      enableColumnFilter: true
    }
    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
    }
    column value #TICKETS {
      label: "TICKETS"
      value: :TICKETS
      enableColumnFilter: true
    }
    column value #PURPOSE_VISIT {
      label: "PURPOSE_VISIT"
      value: :PURPOSE_VISIT
      enableColumnFilter: true
    }
    column value #PURPOSE_VISIT_other {
      label: "PURPOSE_VISIT.98$other"
      value: :PURPOSE_VISIT.98$other
      enableColumnFilter: true
    }
    column value #ARRIVAL_1 {
      label: "ARRIVAL.1"
      value: :ARRIVAL.1
      enableColumnFilter: true
    }
    column value #ARRIVAL_2 {
      label: "ARRIVAL.2"
      value: :ARRIVAL.2
      enableColumnFilter: true
    }
    column value #ARRIVAL_3 {
      label: "ARRIVAL.3"
      value: :ARRIVAL.3
      enableColumnFilter: true
    }
    column value #ARRIVAL_4 {
      label: "ARRIVAL.4"
      value: :ARRIVAL.4
      enableColumnFilter: true
    }
    column value #ARRIVAL_5 {
      label: "ARRIVAL.5"
      value: :ARRIVAL.5
      enableColumnFilter: true
    }
    column value #ARRIVAL_6 {
      label: "ARRIVAL.6"
      value: :ARRIVAL.6
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_attractions {
      label: "SAT_EXPERIENCES.attractions"
      value: :SAT_EXPERIENCES.attractions
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_bars {
      label: "SAT_EXPERIENCES.bars"
      value: :SAT_EXPERIENCES.bars
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_breakfast {
      label: "SAT_EXPERIENCES.breakfast"
      value: :SAT_EXPERIENCES.breakfast
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_bus {
      label: "SAT_EXPERIENCES.bus"
      value: :SAT_EXPERIENCES.bus
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_concierge {
      label: "SAT_EXPERIENCES.concierge"
      value: :SAT_EXPERIENCES.concierge
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_otheramenities {
      label: "SAT_EXPERIENCES.otheramenities"
      value: :SAT_EXPERIENCES.otheramenities
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_premiums {
      label: "SAT_EXPERIENCES.premiums"
      value: :SAT_EXPERIENCES.premiums
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_restaurants {
      label: "SAT_EXPERIENCES.restaurants"
      value: :SAT_EXPERIENCES.restaurants
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_rides {
      label: "SAT_EXPERIENCES.rides"
      value: :SAT_EXPERIENCES.rides
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_shops {
      label: "SAT_EXPERIENCES.shops"
      value: :SAT_EXPERIENCES.shops
      enableColumnFilter: true
    }
    column value #SAT_EXPERIENCES_spa {
      label: "SAT_EXPERIENCES.spa"
      value: :SAT_EXPERIENCES.spa
      enableColumnFilter: true
    }
    column value #ATTRACTIONS_SEEN {
      label: "ATTRACTIONS_SEEN"
      value: :ATTRACTIONS_SEEN
      enableColumnFilter: true
    }
    column value #ATTRACT_INSERT {
      label: "ATTRACT_INSERT"
      value: :ATTRACT_INSERT
      enableColumnFilter: true
    }
    column value #DRILL_ATTRACTION_cleanliness {
      label: "DRILL_ATTRACTION.cleanliness"
      value: :DRILL_ATTRACTION.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_ATTRACTION_quality {
      label: "DRILL_ATTRACTION.quality"
      value: :DRILL_ATTRACTION.quality
      enableColumnFilter: true
    }
    column value #DRILL_ATTRACTION_staff {
      label: "DRILL_ATTRACTION.staff"
      value: :DRILL_ATTRACTION.staff
      enableColumnFilter: true
    }
    column value #DRILL_BUS_cleanarea {
      label: "DRILL_BUS.cleanarea"
      value: :DRILL_BUS.cleanarea
      enableColumnFilter: true
    }
    column value #DRILL_BUS_cleanbus {
      label: "DRILL_BUS.cleanbus"
      value: :DRILL_BUS.cleanbus
      enableColumnFilter: true
    }
    column value #DRILL_BUS_quality {
      label: "DRILL_BUS.quality"
      value: :DRILL_BUS.quality
      enableColumnFilter: true
    }
    column value #DRILL_BUS_staff {
      label: "DRILL_BUS.staff"
      value: :DRILL_BUS.staff
      enableColumnFilter: true
    }
    column value #DRILL_BUS_waitime {
      label: "DRILL_BUS.waitime"
      value: :DRILL_BUS.waitime
      enableColumnFilter: true
    }
    column value #DRILL_SLOTS_avail {
      label: "DRILL_SLOTS.avail"
      value: :DRILL_SLOTS.avail
      enableColumnFilter: true
    }
    column value #DRILL_SLOTS_selection {
      label: "DRILL_SLOTS.selection"
      value: :DRILL_SLOTS.selection
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_avail {
      label: "DRILL_TABLEGAMES.avail"
      value: :DRILL_TABLEGAMES.avail
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_betting {
      label: "DRILL_TABLEGAMES.betting"
      value: :DRILL_TABLEGAMES.betting
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_selection {
      label: "DRILL_TABLEGAMES.selection"
      value: :DRILL_TABLEGAMES.selection
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_staff {
      label: "DRILL_TABLEGAMES.staff"
      value: :DRILL_TABLEGAMES.staff
      enableColumnFilter: true
    }
    column value #DRILL_GAME_DRINK_speed {
      label: "DRILL_GAME_DRINK.speed"
      value: :DRILL_GAME_DRINK.speed
      enableColumnFilter: true
    }
    column value #DRILL_GAME_DRINK_taste {
      label: "DRILL_GAME_DRINK.taste"
      value: :DRILL_GAME_DRINK.taste
      enableColumnFilter: true
    }
    column value #valueColumn_81 {
      label: "DRILL_GAME_DRINK.value"
      value: :DRILL_GAME_DRINK.value
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_accuracy {
      label: "DRILL_LODGING.accuracy"
      value: :DRILL_LODGING.accuracy
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_arrival {
      label: "DRILL_LODGING.arrival"
      value: :DRILL_LODGING.arrival
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_avail {
      label: "DRILL_LODGING.avail"
      value: :DRILL_LODGING.avail
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_cleanliness {
      label: "DRILL_LODGING.cleanliness"
      value: :DRILL_LODGING.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_departure {
      label: "DRILL_LODGING.departure"
      value: :DRILL_LODGING.departure
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_service {
      label: "DRILL_LODGING.service"
      value: :DRILL_LODGING.service
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_staff {
      label: "DRILL_LODGING.staff"
      value: :DRILL_LODGING.staff
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_ac {
      label: "DRILL_ROOM.ac"
      value: :DRILL_ROOM.ac
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathamenities {
      label: "DRILL_ROOM.bathamenities"
      value: :DRILL_ROOM.bathamenities
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathclean {
      label: "DRILL_ROOM.bathclean"
      value: :DRILL_ROOM.bathclean
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathfeatures {
      label: "DRILL_ROOM.bathfeatures"
      value: :DRILL_ROOM.bathfeatures
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bed {
      label: "DRILL_ROOM.bed"
      value: :DRILL_ROOM.bed
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_cleanliness {
      label: "DRILL_ROOM.cleanliness"
      value: :DRILL_ROOM.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_furnishings {
      label: "DRILL_ROOM.furnishings"
      value: :DRILL_ROOM.furnishings
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_quiet {
      label: "DRILL_ROOM.quiet"
      value: :DRILL_ROOM.quiet
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_smell {
      label: "DRILL_ROOM.smell"
      value: :DRILL_ROOM.smell
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_wifi {
      label: "DRILL_ROOM.wifi"
      value: :DRILL_ROOM.wifi
      enableColumnFilter: true
    }
    column value #LODGING_COMMENTS {
      label: "LODGING_COMMENTS"
      value: :LODGING_COMMENTS
      enableColumnFilter: true
    }
    column value #ROOM_COMMENTS {
      label: "ROOM_COMMENTS"
      value: :ROOM_COMMENTS
      enableColumnFilter: true
    }
    column value #RESTAURANT_INSERT {
      label: "RESTAURANT_INSERT"
      value: :RESTAURANT_INSERT
      enableColumnFilter: true
    }
    column value #MEAL_RATED {
      label: "MEAL_RATED"
      value: :MEAL_RATED
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_cleanliness {
      label: "DRILL_RESTAURANT.cleanliness"
      value: :DRILL_RESTAURANT.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_kiosk {
      label: "DRILL_RESTAURANT.kiosk"
      value: :DRILL_RESTAURANT.kiosk
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_quality {
      label: "DRILL_RESTAURANT.quality"
      value: :DRILL_RESTAURANT.quality
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_speed {
      label: "DRILL_RESTAURANT.speed"
      value: :DRILL_RESTAURANT.speed
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_staff {
      label: "DRILL_RESTAURANT.staff"
      value: :DRILL_RESTAURANT.staff
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_value {
      label: "DRILL_RESTAURANT.value"
      value: :DRILL_RESTAURANT.value
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_variety {
      label: "DRILL_RESTAURANT.variety"
      value: :DRILL_RESTAURANT.variety
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_cleanliness {
      label: "DRILL_BUFFET.cleanliness"
      value: :DRILL_BUFFET.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_quality {
      label: "DRILL_BUFFET.quality"
      value: :DRILL_BUFFET.quality
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_stock {
      label: "DRILL_BUFFET.stock"
      value: :DRILL_BUFFET.stock
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_taste {
      label: "DRILL_BUFFET.taste"
      value: :DRILL_BUFFET.taste
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_temperature {
      label: "DRILL_BUFFET.temperature"
      value: :DRILL_BUFFET.temperature
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_value {
      label: "DRILL_BUFFET.value"
      value: :DRILL_BUFFET.value
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_variety {
      label: "DRILL_BUFFET.variety"
      value: :DRILL_BUFFET.variety
      enableColumnFilter: true
    }
    column value #DINING_COMMENT_INSERT {
      label: "DINING_COMMENT_INSERT"
      value: :DINING_COMMENT_INSERT
      enableColumnFilter: true
    }
    column value #RESTAURANT_COMMENTS {
      label: "RESTAURANT_COMMENTS"
      value: :RESTAURANT_COMMENTS
      enableColumnFilter: true
    }
    column value #PREMIUM_PURCHASED {
      label: "PREMIUM_PURCHASED"
      value: :PREMIUM_PURCHASED
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_foodquality {
      label: "DRILL_PREMIUM.foodquality"
      value: :DRILL_PREMIUM.foodquality
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_quality {
      label: "DRILL_PREMIUM.quality"
      value: :DRILL_PREMIUM.quality
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_staff {
      label: "DRILL_PREMIUM.staff"
      value: :DRILL_PREMIUM.staff
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_value {
      label: "DRILL_PREMIUM.value"
      value: :DRILL_PREMIUM.value
      enableColumnFilter: true
    }
    column value #SHOPS_VISITED {
      label: "SHOPS_VISITED"
      value: :SHOPS_VISITED
      enableColumnFilter: true
    }
    column value #SHOPS_INSERT {
      label: "SHOPS_INSERT"
      value: :SHOPS_INSERT
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_merch {
      label: "DRILL_SHOPS.merch"
      value: :DRILL_SHOPS.merch
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_shopsat {
      label: "DRILL_SHOPS.shopsat"
      value: :DRILL_SHOPS.shopsat
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_speed {
      label: "DRILL_SHOPS.speed"
      value: :DRILL_SHOPS.speed
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_staff {
      label: "DRILL_SHOPS.staff"
      value: :DRILL_SHOPS.staff
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_value {
      label: "DRILL_SHOPS.value"
      value: :DRILL_SHOPS.value
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_variety {
      label: "DRILL_SHOPS.variety"
      value: :DRILL_SHOPS.variety
      enableColumnFilter: true
    }
    column value #Problem {
      label: "Problem"
      value: :PROBLEM
      enableColumnFilter: true
    }
    column value #PROB_REPORTED {
      label: "Problem Reported"
      value: :PROB_REPORTED
      enableColumnFilter: true
    }
    column value #RESOLUTION_SAT {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    column value #CONTACT_REQUESTED {
      label: "Contact Requested"
      value: :CONTACT
      enableColumnFilter: true
    }
    column value #CONTACT_PREF {
      label: "Method of Contact"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_name {
      label: "Contact Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_phone {
      label: "Contact Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_email {
      label: "Contact Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #PROBLEM_DETAIL {
      label: "Problem Detail"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #TEAM_REC {
      label: "Team Recognition"
      value: :TEAM_REC
      enableColumnFilter: true
    }
    column value #TEAM_MEMBER {
      label: "Team Member"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #RECOG_DETAIL {
      label: "Team Recognition Detail"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }
    column value #REGION {
      label: "REGION"
      value: :REGION
      enableColumnFilter: true
    }
    column value #GENDER {
      label: "GENDER"
      value: :GENDER
      enableColumnFilter: true
    }
    column value #AGE {
      label: "AGE"
      value: :AGE
      enableColumnFilter: true
    }
    column value #INCOME {
      label: "INCOME"
      value: :INCOME
      enableColumnFilter: true
    }
    column value #UNDER_18_KIDS {
      label: "UNDER_18_KIDS"
      value: :UNDER_18_KIDS
      enableColumnFilter: true
    }
    column value #EDUCATION {
      label: "EDUCATION"
      value: :EDUCATION
      enableColumnFilter: true
    }
    column value #ETHNICITY {
      label: "ETHNICITY"
      value: :ETHNICITY
      enableColumnFilter: true
    }
    column value #COMPANIONS {
      label: "COMPANIONS"
      value: :COMPANIONS
      enableColumnFilter: true
    }
    column value #TOTAL_PARTY {
      label: "TOTAL_PARTY"
      value: :TOTAL_PARTY
      enableColumnFilter: true
    }
    column value #TIME_OF_GAMING_VISIT {
      label: "TIME_OF_GAMING_VISIT"
      value: :TIME_OF_GAMING_VISIT
      enableColumnFilter: true
    }
    column value #WIN_LOSE {
      label: "WIN_LOSE"
      value: :WIN_LOSE
      enableColumnFilter: true
    }
    column value #SPEC_EVENT {
      label: "SPEC_EVENT"
      value: :SPEC_EVENT
      enableColumnFilter: true
    }
    column value #SPEC_EVENT_other {
      label: "SPEC_EVENT.98$other"
      value: :SPEC_EVENT.98$other
      enableColumnFilter: true
    }
    column value #COMPS {
      label: "COMPS"
      value: :COMPS
      enableColumnFilter: true
    }
    column value #COMPS_other {
      label: "COMPS.98$other"
      value: :COMPS.98$other
      enableColumnFilter: true
    }
    column value #REDEMPTION {
      label: "REDEMPTION"
      value: :REDEMPTION
      enableColumnFilter: true
    }
    column value #REDEMPTION_other {
      label: "REDEMPTION.98$other"
      value: :REDEMPTION.98$other
      enableColumnFilter: true
    }
    column value #NO_VISITS {
      label: "NO_VISITS"
      value: :NO_VISITS
      enableColumnFilter: true
    }
    column value #AWARENESS {
      label: "AWARENESS"
      value: :AWARENESS
      enableColumnFilter: true
    }
    column value #KSC_COMPANIONS {
      label: "KSC_COMPANIONS"
      value: :KSC_COMPANIONS
      enableColumnFilter: true
    }
    column value #ACCOMMODATIONS {
      label: "ACCOMMODATIONS"
      value: :ACCOMMODATIONS
      enableColumnFilter: true
    }
    column value #KSC_LOCATION {
      label: "LOCATION"
      value: :LOCATION
      enableColumnFilter: true
    }
    column value #OTHER_ATTRACTIONS {
      label: "OTHER_ATTRACTIONS"
      value: :OTHER_ATTRACTIONS
      enableColumnFilter: true
    }
    column value #NO_VACATIONS {
      label: "NO_VACATIONS"
      value: :NO_VACATIONS
      enableColumnFilter: true
    }


    column value #email {
      label: "email"
      value: :email
      enableColumnFilter: true
    }
    column value #customer_id {
      label: "customer_id"
      value: :customer_id
      enableColumnFilter: true
    }
    column value #player_id {
      label: "player_id"
      value: :player_id
      enableColumnFilter: true
    }
    column value #guest_name {
      label: "guest_name"
      value: :guest_name
      enableColumnFilter: true
    }
    column value #guest_gender {
      label: "guest_gender"
      value: :guest_gender
      enableColumnFilter: true
    }
    column value #customer_state {
      label: "customer_state"
      value: :customer_state
      enableColumnFilter: true
    }
    column value #Postal {
      label: "Postal"
      value: :Postal
      enableColumnFilter: true
    }
    column value #customer_country {
      label: "customer_country"
      value: :customer_country
      enableColumnFilter: true
    }
    column value #customer_city {
      label: "customer_city"
      value: :customer_city
      enableColumnFilter: true
    }
    column value #date_of_birth {
      label: "date_of_birth"
      value: :date_of_birth
      enableColumnFilter: true
    }
    column value #guest_age {
      label: "guest_age"
      value: :guest_age
      enableColumnFilter: true
    }
    column value #TransactionID {
      label: "TransactionID"
      value: :TransactionID
      enableColumnFilter: true
    }
    column value #transaction_time_stamp {
      label: "transaction_time_stamp"
      value: :transaction_time_stamp
      enableColumnFilter: true
    }
    column value #YieldDateTime {
      label: "YieldDateTime"
      value: :YieldDateTime
      enableColumnFilter: true
    }
    column value #CountryName {
      label: "CountryName"
      value: :CountryName
      enableColumnFilter: true
    }
    column value #CompanyID {
      label: "CompanyID"
      value: :CompanyID
      enableColumnFilter: true
    }
    column value #NodeNo {
      label: "NodeNo"
      value: :NodeNo
      enableColumnFilter: true
    }
    column value #SellingPrice {
      label: "SellingPrice"
      value: :SellingPrice
      enableColumnFilter: true
    }
    column value #UseNo {
      label: "UseNo"
      value: :UseNo
      enableColumnFilter: true
    }
    column value #visits {
      label: "visits"
      value: :visits
      enableColumnFilter: true
    }
    column value #minutes_played {
      label: "minutes_played"
      value: :minutes_played
      enableColumnFilter: true
    }
    column value #avgADT {
      label: "avgADT"
      value: :avgADT
      enableColumnFilter: true
    }
    column value #game_pref {
      label: "game_pref"
      value: :game_pref
      enableColumnFilter: true
    }
    column value #rank_description {
      label: "rank_description"
      value: :rank_description
      enableColumnFilter: true
    }
    column value #last_play_date {
      label: "last_play_date"
      value: :last_play_date
      enableColumnFilter: true
    }
    column value #date_enrolled {
      label: "date_enrolled"
      value: :date_enrolled
      enableColumnFilter: true
    }
    column value #total_guest_count {
      label: "total_guest_count"
      value: :total_guest_count
      enableColumnFilter: true
    }
    column value #children_count {
      label: "children_count"
      value: :children_count
      enableColumnFilter: true
    }
    column value #adult_count {
      label: "adult_count"
      value: :adult_count
      enableColumnFilter: true
    }
    column value #reservation_revenue {
      label: "reservation_revenue"
      value: :reservation_revenue
      enableColumnFilter: true
    }
    column value #market_segment_code {
      label: "market_segment_code"
      value: :market_segment_code
      enableColumnFilter: true
    }
    column value #reservation_status {
      label: "reservation_status"
      value: :reservation_status
      enableColumnFilter: true
    }
    column value #room_description {
      label: "room_description"
      value: :room_description
      enableColumnFilter: true
    }
    column value #room_category {
      label: "room_category"
      value: :room_category
      enableColumnFilter: true
    }
    column value #rate_description {
      label: "rate_description"
      value: :rate_description
      enableColumnFilter: true
    }
    column value #departure_date {
      label: "departure_date"
      value: :departure_date
      enableColumnFilter: true
    }
    column value #arrival_date {
      label: "arrival_date"
      value: :arrival_date
      enableColumnFilter: true
    }
    column value #confirm_number {
      label: "confirm_number"
      value: :confirm_number
      enableColumnFilter: true
    }
  } //end widget
  hide: true
  modal: false
} // end page
page #page_GamingResponses {

  label: "Gaming - Response Details"

  widget table #tableWidget {
    label: "Gaming Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start
    rowsPerPage: 100, 500, 1000
    navigateTo: page_Indiv_Survey_Response

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_GamingSurvey()
      label: "Gaming survey Only"
    }

    filter expression {
      value: surveyDataset:filterMeasure_NPSanswered()
      label: "NPS has a value"
    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
    }

    column value #LocationName {
      label: "Location Name"
      value: :LocationName
      enableColumnFilter: true
    }

    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
    }

    column value #RETURN_VISIT {
      label: "Return Visit"
      value: :RETURN_VISIT
      enableColumnFilter: true
    }
    column value #SAT {
      label: "Overall Sat"
      value: :SAT
      enableColumnFilter: true
    }
    column value #GAMING_EXPERIENCES {
      label: "Gaming_Experiences"
      value: :GAMING_EXPERIENCES
      enableColumnFilter: true
    }
    column value #GamingSurveyPath {
      label: "Gaming-Survey Path"
      value: :GamingSurveyPath
      enableColumnFilter: true
    }
    column value #Value {
      label: "Value"
      value: :Value
      enableColumnFilter: true
    }

    column value #SAT_DRIVERS_cleanliness {
      label: "Sat-Cleanliness"
      value: :SAT_DRIVERS.cleanliness
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_safety {
      label: "Sat-Safety"
      value: :SAT_DRIVERS.safety
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_speed {
      label: "Sat-Speed of service"
      value: :SAT_DRIVERS.speed
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_staff {
      label: "Sat-Staff"
      value: :SAT_DRIVERS.staff
      enableColumnFilter: true
    }
    column value #SAT_GAMING_bars {
      label: "Sat-Bars"
      value: :SAT_GAMING.bars
      enableColumnFilter: true
    }
    column value #SAT_GAMING_betting {
      label: "Sat-Betting"
      value: :SAT_GAMING.betting
      enableColumnFilter: true
    }
    column value #SAT_GAMING_buffet {
      label: "Sat-Buffet"
      value: :SAT_GAMING.buffet
      enableColumnFilter: true
    }
    column value #SAT_GAMING_drinks {
      label: "Sat-Drinks"
      value: :SAT_GAMING.drinks
      enableColumnFilter: true
    }
    column value #SAT_GAMING_gaming {
      label: "Sat-Gaming"
      value: :SAT_GAMING.gaming
      enableColumnFilter: true
    }
    column value #SAT_GAMING_lodging {
      label: "Sat-Lodging"
      value: :SAT_GAMING.lodging
      enableColumnFilter: true
    }
    column value #SAT_GAMING_playersclub {
      label: "Sat-Players Club"
      value: :SAT_GAMING.playersclub
      enableColumnFilter: true
    }
    column value #SAT_GAMING_pokerroom {
      label: "Sat-Poker Room"
      value: :SAT_GAMING.pokerroom
      enableColumnFilter: true
    }
    column value #SAT_GAMING_restaurants {
      label: "Sat-Restaurants"
      value: :SAT_GAMING.restaurants
      enableColumnFilter: true
    }
    column value #SAT_GAMING_slots {
      label: "Sat-Slots"
      value: :SAT_GAMING.slots
      enableColumnFilter: true
    }
    column value #SAT_GAMING_tablegames {
      label: "Sat-Table Games"
      value: :SAT_GAMING.tablegames
      enableColumnFilter: true
    }
    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
    }
    column value #DRILL_SLOTS_avail {
      label: "Slots-Availability"
      value: :DRILL_SLOTS.avail
      enableColumnFilter: true
    }
    column value #DRILL_SLOTS_selection {
      label: "Slots-Selection"
      value: :DRILL_SLOTS.selection
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_avail {
      label: "Table Games-Availability"
      value: :DRILL_TABLEGAMES.avail
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_betting {
      label: "Table Games-Betting"
      value: :DRILL_TABLEGAMES.betting
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_selection {
      label: "Table Games-Selection"
      value: :DRILL_TABLEGAMES.selection
      enableColumnFilter: true
    }
    column value #DRILL_TABLEGAMES_staff {
      label: "Table Games-Staff"
      value: :DRILL_TABLEGAMES.staff
      enableColumnFilter: true
    }
    column value #DRILL_GAME_DRINK_speed {
      label: "Drinks-Speed of servce"
      value: :DRILL_GAME_DRINK.speed
      enableColumnFilter: true
    }
    column value #DRILL_GAME_DRINK_taste {
      label: "Drinks-Taste"
      value: :DRILL_GAME_DRINK.taste
      enableColumnFilter: true
    }
    column value #valueColumn_81 {
      label: "Drinks-Value"
      value: :DRILL_GAME_DRINK.value
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_accuracy {
      label: "Lodging-Reservation accuracy"
      value: :DRILL_LODGING.accuracy
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_arrival {
      label: "Lodging-Arrival experience"
      value: :DRILL_LODGING.arrival
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_avail {
      label: "Lodging-Staff availability"
      value: :DRILL_LODGING.avail
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_cleanliness {
      label: "Lodging-Cleanliness"
      value: :DRILL_LODGING.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_departure {
      label: "Lodging-Departure experience"
      value: :DRILL_LODGING.departure
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_service {
      label: "Lodging-Service"
      value: :DRILL_LODGING.service
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_staff {
      label: "Lodging-Staff"
      value: :DRILL_LODGING.staff
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_ac {
      label: "Room-A/C-Heating"
      value: :DRILL_ROOM.ac
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathamenities {
      label: "Room-Bath Amenities"
      value: :DRILL_ROOM.bathamenities
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathclean {
      label: "Room-Clean bath"
      value: :DRILL_ROOM.bathclean
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathfeatures {
      label: "Room-Bath features"
      value: :DRILL_ROOM.bathfeatures
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bed {
      label: "Room-Bed"
      value: :DRILL_ROOM.bed
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_cleanliness {
      label: "Room-Cleanliness"
      value: :DRILL_ROOM.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_furnishings {
      label: "Room-Furnishings"
      value: :DRILL_ROOM.furnishings
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_quiet {
      label: "Room-Quiet"
      value: :DRILL_ROOM.quiet
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_smell {
      label: "Room-Smell"
      value: :DRILL_ROOM.smell
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_wifi {
      label: "Room-Wifi"
      value: :DRILL_ROOM.wifi
      enableColumnFilter: true
    }
    column value #LODGING_COMMENTS {
      label: "Lodging Comments"
      value: :LODGING_COMMENTS
      enableColumnFilter: true
    }

    column value #RESTAURANT_INSERT {
      label: "RESTAURANT INSERT"
      value: :RESTAURANT_INSERT
      enableColumnFilter: true
    }
    column value #MEAL_RATED {
      label: "Meal Rated"
      value: :MEAL_RATED
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_cleanliness {
      label: "Restaurant-Cleanliness"
      value: :DRILL_RESTAURANT.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_kiosk {
      label: "Restaurant-Kiosk"
      value: :DRILL_RESTAURANT.kiosk
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_quality {
      label: "Restaurant-Quality of food/bev"
      value: :DRILL_RESTAURANT.quality
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_speed {
      label: "Restaurant-Speed of service"
      value: :DRILL_RESTAURANT.speed
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_staff {
      label: "Restaurant-Staff"
      value: :DRILL_RESTAURANT.staff
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_value {
      label: "Restaurant-Value"
      value: :DRILL_RESTAURANT.value
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_variety {
      label: "Restaurant-Variety"
      value: :DRILL_RESTAURANT.variety
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_cleanliness {
      label: "Buffet-Cleanliness"
      value: :DRILL_BUFFET.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_quality {
      label: "Buffet-Quality"
      value: :DRILL_BUFFET.quality
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_stock {
      label: "Buffet-Well-stocked"
      value: :DRILL_BUFFET.stock
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_taste {
      label: "Buffet-Taste"
      value: :DRILL_BUFFET.taste
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_temperature {
      label: "Buffet-Temperature"
      value: :DRILL_BUFFET.temperature
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_value {
      label: "Buffet-Value"
      value: :DRILL_BUFFET.value
      enableColumnFilter: true
    }
    column value #DRILL_BUFFET_variety {
      label: "Buffet-Variety"
      value: :DRILL_BUFFET.variety
      enableColumnFilter: true
    }

    column value #RESTAURANT_COMMENTS {
      label: "Restaurant Comments"
      value: :RESTAURANT_COMMENTS
      enableColumnFilter: true
    }

    column value #Problem {
      label: "Problem"
      value: :PROBLEM
      enableColumnFilter: true
    }
    column value #PROB_REPORTED {
      label: "Problem Reported"
      value: :PROB_REPORTED
      enableColumnFilter: true
    }
    column value #RESOLUTION_SAT {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    column value #CONTACT_REQUESTED {
      label: "Contact Requested"
      value: :CONTACT
      enableColumnFilter: true
    }
    column value #CONTACT_PREF {
      label: "Method of Contact"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_name {
      label: "Contact Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_phone {
      label: "Contact Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_email {
      label: "Contact Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #PROBLEM_DETAIL {
      label: "Problem Detail"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #TEAM_REC {
      label: "Team Recognition"
      value: :TEAM_REC
      enableColumnFilter: true
    }
    column value #TEAM_MEMBER {
      label: "Team Member"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #RECOG_DETAIL {
      label: "Team Recognition Detail"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }
  //begin demos
    column value #REGION {
      label: "REGION"
      value: :REGION
      enableColumnFilter: true
    }
    column value #GENDER {
      label: "GENDER"
      value: :GENDER
      enableColumnFilter: true
    }
    column value #AGE {
      label: "AGE"
      value: :AGE
      enableColumnFilter: true
    }
    column value #INCOME {
      label: "INCOME"
      value: :INCOME
      enableColumnFilter: true
    }
    column value #UNDER_18_KIDS {
      label: "NUM CHILDREN"
      value: :UNDER_18_KIDS
      enableColumnFilter: true
    }
    column value #EDUCATION {
      label: "EDUCATION"
      value: :EDUCATION
      enableColumnFilter: true
    }
    column value #ETHNICITY {
      label: "ETHNICITY"
      value: :ETHNICITY
      enableColumnFilter: true
    }
    column value #COMPANIONS {
      label: "COMPANIONS"
      value: :COMPANIONS
      enableColumnFilter: true
    }
    column value #TOTAL_PARTY {
      label: "NUM IN TOTAL PARTY"
      value: :TOTAL_PARTY
      enableColumnFilter: true
    }
    column value #TIME_OF_GAMING_VISIT {
      label: "TIME OF GAMING VISIT"
      value: :TIME_OF_GAMING_VISIT
      enableColumnFilter: true
    }
    column value #WIN_LOSE {
      label: "WIN OR LOSE"
      value: :WIN_LOSE
      enableColumnFilter: true
    }
    column value #SPEC_EVENT {
      label: "SPECIAL EVENT"
      value: :SPEC_EVENT
      enableColumnFilter: true
    }
    column value #SPEC_EVENT_other {
      label: "SPECIAL EVENT-OTHER"
      value: :SPEC_EVENT.98$other
      enableColumnFilter: true
    }
    column value #COMPS {
      label: "COMPS"
      value: :COMPS
      enableColumnFilter: true
    }
    column value #COMPS_other {
      label: "COMPS-OTHER"
      value: :COMPS.98$other
      enableColumnFilter: true
    }
    column value #REDEMPTION {
      label: "REDEMPTION"
      value: :REDEMPTION
      enableColumnFilter: true
    }
    column value #REDEMPTION_other {
      label: "REDEMPTION-OTHER"
      value: :REDEMPTION.98$other
      enableColumnFilter: true
    }
//begin background info
    column value #email {
      label: "email"
      value: :email
      enableColumnFilter: true
    }
    column value #customer_id {
      label: "Customer id"
      value: :customer_id
      enableColumnFilter: true
    }
    column value #player_id {
      label: "Player id"
      value: :player_id
      enableColumnFilter: true
    }
    column value #guest_name {
      label: "Guest name"
      value: :guest_name
      enableColumnFilter: true
    }
    column value #guest_gender {
      label: "Guest gender"
      value: :guest_gender
      enableColumnFilter: true
    }
    column value #customer_state {
      label: "Customer state"
      value: :customer_state
      enableColumnFilter: true
    }
    column value #Postal {
      label: "Customer postal"
      value: :Postal
      enableColumnFilter: true
    }
    column value #customer_country {
      label: "Customer country"
      value: :customer_country
      enableColumnFilter: true
    }
    column value #customer_city {
      label: "Customer city"
      value: :customer_city
      enableColumnFilter: true
    }
    column date #date_of_birth {
      label: "Date of birth"
      value: :date_of_birth
      enableColumnFilter: true
    }
    column value #guest_age {
      label: "Guest age"
      value: :guest_age
      enableColumnFilter: true
    }
    column value #TransactionID {
      label: "Transaction ID"
      value: :TransactionID
      enableColumnFilter: true
    }
    column value #transaction_time_stamp {
      label: "Transaction date"
      value: :transaction_time_stamp
      enableColumnFilter: true
    }
    column value #visits {
      label: "Num visits"
      value: :visits
      enableColumnFilter: true
    }
    column value #minutes_played {
      label: "Minutes played"
      value: :minutes_played
      enableColumnFilter: true
    }
    column value #avgADT {
      label: "Avg ADT"
      value: :avgADT
      enableColumnFilter: true
    }
    column value #game_pref {
      label: "Game pref"
      value: :game_pref
      enableColumnFilter: true
    }
    column value #rank_description {
      label: "Loyalty tier"
      value: :rank_description
      enableColumnFilter: true
    }
    column date #last_play_date {
      label: "Last play date"
      value: :last_play_date
      enableColumnFilter: true
    }
    column date #date_enrolled {
      label: "Date enrolled"
      value: :date_enrolled
      enableColumnFilter: true
    }
    column value #total_guest_count {
      label: "Total guest count"
      value: :total_guest_count
      enableColumnFilter: true
    }
    column value #children_count {
      label: "Children count"
      value: :children_count
      enableColumnFilter: true
    }
    column value #adult_count {
      label: "Adult count"
      value: :adult_count
      enableColumnFilter: true
    }
    column value #reservation_revenue {
      label: "Reservation revenue"
      value: :reservation_revenue
      enableColumnFilter: true
    }
    column value #market_segment_code {
      label: "Market segment code"
      value: :market_segment_code
      enableColumnFilter: true
    }
    column value #reservation_status {
      label: "Reservation status"
      value: :reservation_status
      enableColumnFilter: true
    }
    column value #room_description {
      label: "Room description"
      value: :room_description
      enableColumnFilter: true
    }
    column value #room_category {
      label: "Room category"
      value: :room_category
      enableColumnFilter: true
    }
    column value #rate_description {
      label: "Rate description"
      value: :rate_description
      enableColumnFilter: true
    }
    column date #departure_date {
      label: "Departure date"
      value: :departure_date
      enableColumnFilter: true
    }
    column date #arrival_date {
      label: "Arrival date"
      value: :arrival_date
      enableColumnFilter: true
    }
    column value #confirm_number {
      label: "Confirm number"
      value: :confirm_number
      enableColumnFilter: true
    }
  } //end widget
  hide: false
  modal: true
} // end page
page #page_SouthlandSegmentationResponses {

  label: "Southland Gaming Segmentation Response Details"

  widget table #tableWidget {
    label: "Southland Casino Hotel Personas Segmentation Drilldown"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start
    rowsPerPage: 100, 500, 1000
    navigateTo: page_Indiv_Survey_Response

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_GamingSurvey()
      label: "Gaming survey Only"
    }

    filter expression {
      value: surveyDataset:filterMeasure_NPSanswered()
      label: "NPS has a value"
    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
      align: center
    }

    column value #LocationName {
      label: "Location Name"
      value: :LocationName
      enableColumnFilter: true
      align: center
    }

    column value #SOUTHLAND_SEGMENTATION_assign {
      label: "Southland Persona"
      value: :Southland_Gaming_Seg_assign
      enableColumnFilter: true
      align: center
    }

    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
      align: center
    }

    column value #SAT {
      label: "Overall Sat"
      value: :SAT
      enableColumnFilter: true
      align: center
    }

    column value #SOUTHLAND_SEGMENTATION_fun {
      label: "Reason to visit-Fun Experience"
      value: :GAMING_SEGMENTATION.funexperience
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_winagain {
      label: "Reason to visit-Win Again"
      value: :GAMING_SEGMENTATION.winagain
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_relax {
      label: "Reason to visit-Relax"
      value: :GAMING_SEGMENTATION.relax
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_entertain {
      label: "Reason to visit-Entertain others"
      value: :GAMING_SEGMENTATION.entertain
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_lifechanging {
      label: "Reason to visit-Life Changing"
      value: :GAMING_SEGMENTATION.lifechanging
      enableColumnFilter: true
      align: center
    }

    column value #SOUTHLAND_SEGMENTATION_overnightstay {
      label: "Reason to visit-Vacation"
      value: :GAMING_SEGMENTATION.overnightstay
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_skills {
      label: "Reason to visit-Skills"
      value: :GAMING_SEGMENTATION.skills
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_funalone {
      label: "Reason to visit-Fun Alone"
      value: :GAMING_SEGMENTATION.funalone
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_tobesurprised {
      label: "Reason to visit-To Be Surprised"
      value: :GAMING_SEGMENTATION.tobesurprised
      enableColumnFilter: true
      align: center
    }
    column value #SOUTHLAND_SEGMENTATION_treatmyself {
      label: "Reason to visit-Treat Myself"
      value: :GAMING_SEGMENTATION.treatmyself
      enableColumnFilter: true
      align: center
    }

    column value #REGION {
      label: "REGION"
      value: :REGION
      enableColumnFilter: true
    }
    column value #GENDER {
      label: "GENDER"
      value: :GENDER
      enableColumnFilter: true
    }
    column value #AGE {
      label: "AGE"
      value: :AGE
      enableColumnFilter: true
    }
    column value #INCOME {
      label: "INCOME"
      value: :INCOME
      enableColumnFilter: true
    }
    column value #UNDER_18_KIDS {
      label: "NUM CHILDREN"
      value: :UNDER_18_KIDS
      enableColumnFilter: true
    }
    column value #EDUCATION {
      label: "EDUCATION"
      value: :EDUCATION
      enableColumnFilter: true
    }
    column value #ETHNICITY {
      label: "ETHNICITY"
      value: :ETHNICITY
      enableColumnFilter: true
    }
    column value #COMPANIONS {
      label: "COMPANIONS"
      value: :COMPANIONS
      enableColumnFilter: true
    }
    column value #TOTAL_PARTY {
      label: "NUM IN TOTAL PARTY"
      value: :TOTAL_PARTY
      enableColumnFilter: true
    }
    column value #TIME_OF_GAMING_VISIT {
      label: "TIME OF GAMING VISIT"
      value: :TIME_OF_GAMING_VISIT
      enableColumnFilter: true
    }
    column value #WIN_LOSE {
      label: "WIN OR LOSE"
      value: :WIN_LOSE
      enableColumnFilter: true
    }
    column value #SPEC_EVENT {
      label: "SPECIAL EVENT"
      value: :SPEC_EVENT
      enableColumnFilter: true
    }
    column value #SPEC_EVENT_other {
      label: "SPECIAL EVENT-OTHER"
      value: :SPEC_EVENT.98$other
      enableColumnFilter: true
    }
    column value #COMPS {
      label: "COMPS"
      value: :COMPS
      enableColumnFilter: true
    }
    column value #COMPS_other {
      label: "COMPS-OTHER"
      value: :COMPS.98$other
      enableColumnFilter: true
    }
    column value #REDEMPTION {
      label: "REDEMPTION"
      value: :REDEMPTION
      enableColumnFilter: true
    }
    column value #REDEMPTION_other {
      label: "REDEMPTION-OTHER"
      value: :REDEMPTION.98$other
      enableColumnFilter: true
    }

    column value #email {
      label: "email"
      value: :email
      enableColumnFilter: true
    }
    column value #customer_id {
      label: "Customer id"
      value: :customer_id
      enableColumnFilter: true
    }
    column value #player_id {
      label: "Player id"
      value: :player_id
      enableColumnFilter: true
    }
    column value #guest_name {
      label: "Guest name"
      value: :guest_name
      enableColumnFilter: true
    }
    column value #guest_gender {
      label: "Guest gender"
      value: :guest_gender
      enableColumnFilter: true
    }
    column value #customer_state {
      label: "Customer state"
      value: :customer_state
      enableColumnFilter: true
    }
    column value #Postal {
      label: "Customer postal"
      value: :Postal
      enableColumnFilter: true
    }
    column value #customer_country {
      label: "Customer country"
      value: :customer_country
      enableColumnFilter: true
    }
    column value #customer_city {
      label: "Customer city"
      value: :customer_city
      enableColumnFilter: true
    }
    column date #date_of_birth {
      label: "Date of birth"
      value: :date_of_birth
      enableColumnFilter: true
    }
    column value #guest_age {
      label: "Guest age"
      value: :guest_age
      enableColumnFilter: true
    }
    column value #TransactionID {
      label: "Transaction ID"
      value: :TransactionID
      enableColumnFilter: true
    }
    column value #transaction_time_stamp {
      label: "Transaction date"
      value: :transaction_time_stamp
      enableColumnFilter: true
    }
    column value #visits {
      label: "Num visits"
      value: :visits
      enableColumnFilter: true
    }
    column value #minutes_played {
      label: "Minutes played"
      value: :minutes_played
      enableColumnFilter: true
    }
    column value #avgADT {
      label: "Avg ADT"
      value: :avgADT
      enableColumnFilter: true
    }
    column value #game_pref {
      label: "Game pref"
      value: :game_pref
      enableColumnFilter: true
    }
    column value #rank_description {
      label: "Loyalty tier"
      value: :rank_description
      enableColumnFilter: true
    }
    column date #last_play_date {
      label: "Last play date"
      value: :last_play_date
      enableColumnFilter: true
    }
    column date #date_enrolled {
      label: "Date enrolled"
      value: :date_enrolled
      enableColumnFilter: true
    }
    column value #total_guest_count {
      label: "Total guest count"
      value: :total_guest_count
      enableColumnFilter: true
    }
    column value #children_count {
      label: "Children count"
      value: :children_count
      enableColumnFilter: true
    }
    column value #adult_count {
      label: "Adult count"
      value: :adult_count
      enableColumnFilter: true
    }
    column value #reservation_revenue {
      label: "Reservation revenue"
      value: :reservation_revenue
      enableColumnFilter: true
    }
    column value #market_segment_code {
      label: "Market segment code"
      value: :market_segment_code
      enableColumnFilter: true
    }
    column value #reservation_status {
      label: "Reservation status"
      value: :reservation_status
      enableColumnFilter: true
    }
    column value #room_description {
      label: "Room description"
      value: :room_description
      enableColumnFilter: true
    }
    column value #room_category {
      label: "Room category"
      value: :room_category
      enableColumnFilter: true
    }
    column value #rate_description {
      label: "Rate description"
      value: :rate_description
      enableColumnFilter: true
    }
    column date #departure_date {
      label: "Departure date"
      value: :departure_date
      enableColumnFilter: true
    }
    column date #arrival_date {
      label: "Arrival date"
      value: :arrival_date
      enableColumnFilter: true
    }
    column value #confirm_number {
      label: "Confirm number"
      value: :confirm_number
      enableColumnFilter: true
    }
  } //end widget
  hide: false
  modal: true
  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_Southland_Gaming_Segs()
    label: "Southland Segments"
  }
} // end page
page #page_LodgingResponses {

  label: "Lodging - Response Details"

  hide: false
  modal: true

  widget table #tableWidget {
    label: "Lodging Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_LodgingSurvey()
      label: "Lodging survey Only"
    }

    filter expression {
      value: surveyDataset:filterMeasure_NPSanswered()
      label: "NPS has a value"
    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
    }

    column value #LocationName {
      label: "Location Name"
      value: :LocationName
      enableColumnFilter: true
    }

    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
    }


    column value #SAT {
      label: "Overall Satisfaction"
      value: :SAT
      enableColumnFilter: true
    }

    column value #Value {
      label: "Value"
      value: :Value
      enableColumnFilter: true
    }


    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
    }

    column value #EXPERIENCES {
      label: "EXPERIENCES"
      value: :EXPERIENCES
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_lodging {
      label: "Sat-Lodging"
      value: :SAT_EXPERIENCES.lodging
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_restaurants {
      label: "Sat-Restaurants"
      value: :SAT_EXPERIENCES.restaurants
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_breakfast {
      label: "Sat-Breakfast"
      value: :SAT_EXPERIENCES.breakfast
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_bars {
      label: "Sat-Bars"
      value: :SAT_EXPERIENCES.bars
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_shops {
      label: "SAT_EXPERIENCES.shops"
      value: :SAT_EXPERIENCES.shops
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_concierge {
      label: "Sat-Concierge"
      value: :SAT_EXPERIENCES.concierge
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_spa {
      label: "Sat-Spa"
      value: :SAT_EXPERIENCES.spa
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_otheramenities {
      label: "Sat-Other amenities"
      value: :SAT_EXPERIENCES.otheramenities
      enableColumnFilter: true
    }


    column value #DRILL_LODGING_accuracy {
      label: "Lodging-Accuracy"
      value: :DRILL_LODGING.accuracy
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_arrival {
      label: "Lodging-Arrival"
      value: :DRILL_LODGING.arrival
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_avail {
      label: "Lodging-Avail"
      value: :DRILL_LODGING.avail
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_cleanliness {
      label: "Lodging-Cleanliness"
      value: :DRILL_LODGING.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_departure {
      label: "Lodging-Departure"
      value: :DRILL_LODGING.departure
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_service {
      label: "Lodging-Service"
      value: :DRILL_LODGING.service
      enableColumnFilter: true
    }
    column value #DRILL_LODGING_staff {
      label: "Lodging-Staff"
      value: :DRILL_LODGING.staff
      enableColumnFilter: true
    }

    column value #LODGING_COMMENTS {
      label: "Lodging-Comments"
      value: :LODGING_COMMENTS
      enableColumnFilter: true
    }

    column value #DRILL_ROOM_ac {
      label: "Room-A/C"
      value: :DRILL_ROOM.ac
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathamenities {
      label: "Room-Bath Amenities"
      value: :DRILL_ROOM.bathamenities
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathclean {
      label: "Room-Bath Clean"
      value: :DRILL_ROOM.bathclean
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bathfeatures {
      label: "Room-Bath Features"
      value: :DRILL_ROOM.bathfeatures
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_bed {
      label: "Room-Bed"
      value: :DRILL_ROOM.bed
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_cleanliness {
      label: "Room-Cleanliness"
      value: :DRILL_ROOM.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_furnishings {
      label: "Room-Furnishings"
      value: :DRILL_ROOM.furnishings
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_quiet {
      label: "Room-Quiet"
      value: :DRILL_ROOM.quiet
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_smell {
      label: "Room-Smell"
      value: :DRILL_ROOM.smell
      enableColumnFilter: true
    }
    column value #DRILL_ROOM_wifi {
      label: "Room-Wifi"
      value: :DRILL_ROOM.wifi
      enableColumnFilter: true
    }

    column value #ROOM_COMMENTS {
      label: "Room-Comments"
      value: :ROOM_COMMENTS
      enableColumnFilter: true
    }
    column value #RESTAURANT_INSERT {
      label: "Restaurant Rated"
      value: :RESTAURANT_INSERT_TEXT
      enableColumnFilter: true
    }
    column value #MEAL_RATED {
      label: "Meal Rated"
      value: :MEAL_RATED
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_cleanliness {
      label: "Restaurant-Cleanliness"
      value: :DRILL_RESTAURANT.cleanliness
      enableColumnFilter: true
    }

    column value #DRILL_RESTAURANT_quality {
      label: "Restaurant-Quality"
      value: :DRILL_RESTAURANT.quality
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_speed {
      label: "Restaurant-Speed"
      value: :DRILL_RESTAURANT.speed
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_staff {
      label: "Restaurant-Staff"
      value: :DRILL_RESTAURANT.staff
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_value {
      label: "Restaurant-Value"
      value: :DRILL_RESTAURANT.value
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_variety {
      label: "Restaurant-Variety"
      value: :DRILL_RESTAURANT.variety
      enableColumnFilter: true
    }

    column value #RESTAURANT_COMMENTS {
      label: "Restaurant-Comments"
      value: :RESTAURANT_COMMENTS
      enableColumnFilter: true
    }

    column value #Problem {
      label: "Problem"
      value: :PROBLEM
      enableColumnFilter: true
    }
    column value #PROB_REPORTED {
      label: "Problem Reported"
      value: :PROB_REPORTED
      enableColumnFilter: true
    }
    column value #RESOLUTION_SAT {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    column value #CONTACT_REQUESTED {
      label: "Contact Requested"
      value: :CONTACT
      enableColumnFilter: true
    }
    column value #CONTACT_PREF {
      label: "Method of Contact"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_name {
      label: "Contact Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_phone {
      label: "Contact Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_email {
      label: "Contact Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #PROBLEM_DETAIL {
      label: "Problem Detail"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #TEAM_REC {
      label: "Team Recognition"
      value: :TEAM_REC
      enableColumnFilter: true
    }
    column value #TEAM_MEMBER {
      label: "Team Member"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #RECOG_DETAIL {
      label: "Team Recognition Detail"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }
    column value #REGION {
      label: "REGION"
      value: :REGION
      enableColumnFilter: true
    }
    column value #GENDER {
      label: "GENDER"
      value: :GENDER
      enableColumnFilter: true
    }
    column value #AGE {
      label: "AGE"
      value: :AGE
      enableColumnFilter: true
    }
    column value #INCOME {
      label: "INCOME"
      value: :INCOME
      enableColumnFilter: true
    }
    column value #UNDER_18_KIDS {
      label: "UNDER 18-KIDS"
      value: :UNDER_18_KIDS
      enableColumnFilter: true
    }
    column value #EDUCATION {
      label: "EDUCATION"
      value: :EDUCATION
      enableColumnFilter: true
    }
    column value #ETHNICITY {
      label: "ETHNICITY"
      value: :ETHNICITY
      enableColumnFilter: true
    }
    column value #NO_VISITS {
      label: "NUM VISITS"
      value: :NO_VISITS
      enableColumnFilter: true
    }
    column value #COMPANIONS {
      label: "COMPANIONS"
      value: :COMPANIONS
      enableColumnFilter: true
    }
    column value #NO_VACATIONS {
      label: "NUM VACATIONS"
      value: :NO_VACATIONS
      enableColumnFilter: true
    }

    column value #email {
      label: "email"
      value: :email
      enableColumnFilter: true
    }
    column value #customer_id {
      label: "customer id"
      value: :customer_id
      enableColumnFilter: true
    }

    column value #guest_name {
      label: "guest name"
      value: :guest_name
      enableColumnFilter: true
    }
    column value #guest_gender {
      label: "guest gender"
      value: :guest_gender
      enableColumnFilter: true
    }
    column value #customer_state {
      label: "customer state"
      value: :customer_state
      enableColumnFilter: true
    }
    column value #Postal {
      label: "Postal"
      value: :Postal
      enableColumnFilter: true
    }
    column value #customer_country {
      label: "customer country"
      value: :customer_country
      enableColumnFilter: true
    }
    column value #customer_city {
      label: "customer city"
      value: :customer_city
      enableColumnFilter: true
    }
    column value #transaction_time_stamp {
      label: "transaction time stamp"
      value: :transaction_time_stamp
      enableColumnFilter: true
    }
    column value #total_guest_count {
      label: "total guest count"
      value: :total_guest_count
      enableColumnFilter: true
    }
    column value #children_count {
      label: "children count"
      value: :children_count
      enableColumnFilter: true
    }
    column value #adult_count {
      label: "adult count"
      value: :adult_count
      enableColumnFilter: true
    }
    column value #reservation_revenue {
      label: "reservation revenue"
      value: :reservation_revenue
      enableColumnFilter: true
    }
    column value #market_segment_code {
      label: "market segment code"
      value: :market_segment_code
      enableColumnFilter: true
    }
    column value #reservation_status {
      label: "reservation status"
      value: :reservation_status
      enableColumnFilter: true
    }
    column value #room_description {
      label: "room description"
      value: :room_description
      enableColumnFilter: true
    }
    column value #room_category {
      label: "room category"
      value: :room_category
      enableColumnFilter: true
    }
    column value #rate_description {
      label: "rate description"
      value: :rate_description
      enableColumnFilter: true
    }
    column date #departure_date {
      label: "departure date"
      value: :departure_date
      enableColumnFilter: true
    }
    column date #arrival_date {
      label: "arrival date"
      value: :arrival_date
      enableColumnFilter: true
    }
    column value #confirm_number {
      label: "confirm number"
      value: :confirm_number
      enableColumnFilter: true
    }
    navigateTo: page_Indiv_Survey_Response
  } //end widget
} // end page
page #page_ToursResponses {

  label: "Tours - Response Details"

  hide: false
  modal: true

  widget table #tableWidget {
    label: "Tours and Activities Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_ToursSurvey()
      label: "Lodging survey Only"
    }

    filter expression {
      value: surveyDataset:filterMeasure_NPSanswered()
      label: "NPS has a value"
    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
    }

    column value #LocationName {
      label: "Location Name"
      value: :LocationName
      enableColumnFilter: true
    }


    column value #TourActivityName {
      label: "Tour Activity Name"
      value: :TourActivityName
      enableColumnFilter: true
    }

    column date #TourVisitDate {
      label: "Tour Visit Date"
      value: :TourVisitDate
      enableColumnFilter: true
    }

    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
    }

    column value #SAT {
      label: "Overall Satisfaction"
      value: :SAT
      enableColumnFilter: true
    }

    column value #Value {
      label: "Value"
      value: :Value
      enableColumnFilter: true
    }

    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
    }

    column value #BOOKING_METHOD {
      label: "Booking Method"
      value: :BOOKING_METHOD
      enableColumnFilter: true
    }

    column value #DRILL_BOOKING_SAT {
      label: "Booking-Sat"
      value: :DRILL_BOOKING.bookingsat
      enableColumnFilter: true
    }

    column value #DRILL_BOOKING_availability {
      label: "Booking-Availability"
      value: :DRILL_BOOKING.avail
      enableColumnFilter: true
    }

    column value #DRILL_BOOKING_info {
      label: "Booking-Info"
      value: :DRILL_BOOKING.info
      enableColumnFilter: true
    }

    column value #DRILL_BOOKING_communication {
      label: "Booking-Communication"
      value: :DRILL_BOOKING.communication
      enableColumnFilter: true
    }

    column value #BOOKING_COMMENTS {
      label: "Booking Comments"
      value: :BOOKING_COMMENTS
      enableColumnFilter: true
    }

    column value #DRILL_TOURS_avail {
      label: "Tours-Availability"
      value: :DRILL_TOURS.avail
      enableColumnFilter: true
    }

    column value #DRILL_TOURS_staff {
      label: "Tours-Staff"
      value: :DRILL_TOURS.staff
      enableColumnFilter: true
    }

    column value #DRILL_TOURS_knowledge {
      label: "Tours-Availability"
      value: :DRILL_TOURS.knowledge
      enableColumnFilter: true
    }

    column value #DRILL_TOURS_equipment {
      label: "Tours-Equipment"
      value: :DRILL_TOURS.equipment
      enableColumnFilter: true
    }

    column value #TOURS_COMMENTS {
      label: "Tours Comments"
      value: :TOURS_COMMENTS
      enableColumnFilter: true
    }

    column value #TOURS_ELEMENTS_guidesat {
      label: "Tour Guide-Sat"
      value: :TOURS_ELEMENTS.guidesat
      enableColumnFilter: true
    }

    column value #TOURS_ELEMENTS_knowledge {
      label: "Tour Guide-Knowledge"
      value: :TOURS_ELEMENTS.knowledge
      enableColumnFilter: true
    }

    column value #TOURS_ELEMENTS_toursafety {
      label: "Tour-Safety"
      value: :TOURS_ELEMENTS.toursafety
      enableColumnFilter: true
    }
    column value #TOURS_ELEMENTS_sitesat {
      label: "Tour Sites-Sat"
      value: :TOURS_ELEMENTS.sitesat
      enableColumnFilter: true
    }
    column value #TOURS_ELEMENTS_cleanbus {
      label: "Tour-Clean Vehicle"
      value: :TOURS_ELEMENTS.cleanbus
      enableColumnFilter: true
    }
    column value #TOURS_ELEMENTS_lunch {
      label: "Tour-Lunch"
      value: :TOURS_ELEMENTS.lunch
      enableColumnFilter: true
    }

    column value #ELEMENTS_COMMENT {
      label: "Elements Comments"
      value: :ELEMENTS_COMMENT
      enableColumnFilter: true
    }

    column value #Problem {
      label: "Problem"
      value: :PROBLEM
      enableColumnFilter: true
    }
    column value #PROB_REPORTED {
      label: "Problem Reported"
      value: :PROB_REPORTED
      enableColumnFilter: true
    }
    column value #RESOLUTION_SAT {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    column value #CONTACT_REQUESTED {
      label: "Contact Requested"
      value: :CONTACT
      enableColumnFilter: true
    }
    column value #CONTACT_PREF {
      label: "Method of Contact"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_name {
      label: "Contact Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_phone {
      label: "Contact Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_email {
      label: "Contact Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #PROBLEM_DETAIL {
      label: "Problem Detail"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #TEAM_REC {
      label: "Team Recognition"
      value: :TEAM_REC
      enableColumnFilter: true
    }
    column value #TEAM_MEMBER {
      label: "Team Member"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #RECOG_DETAIL {
      label: "Team Recognition Detail"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }
    column value #REGION {
      label: "REGION"
      value: :REGION
      enableColumnFilter: true
    }
    column value #GENDER {
      label: "GENDER"
      value: :GENDER
      enableColumnFilter: true
    }
    column value #AGE {
      label: "AGE"
      value: :AGE
      enableColumnFilter: true
    }
    column value #INCOME {
      label: "INCOME"
      value: :INCOME
      enableColumnFilter: true
    }
    column value #UNDER_18_KIDS {
      label: "UNDER 18-KIDS"
      value: :UNDER_18_KIDS
      enableColumnFilter: true
    }
    column value #EDUCATION {
      label: "EDUCATION"
      value: :EDUCATION
      enableColumnFilter: true
    }
    column value #ETHNICITY {
      label: "ETHNICITY"
      value: :ETHNICITY
      enableColumnFilter: true
    }

    column value #NO_VISITS {
      label: "NUM VISITS"
      value: :NO_VISITS
      enableColumnFilter: true
    }

    column value #ADVANCE_BOOKING {
      label: "ADVANCE BOOKING"
      value: :ADVANCE_BOOKING
      enableColumnFilter: true
    }

    column value #COMPANIONS {
      label: "COMPANIONS"
      value: :COMPANIONS
      enableColumnFilter: true
    }
    column value #NO_VACATIONS {
      label: "NUM VACATIONS"
      value: :NO_VACATIONS
      enableColumnFilter: true
    }

    column value #email {
      label: "email"
      value: :email
      enableColumnFilter: true
    }
    column value #customer_id {
      label: "customer id"
      value: :CustomerID
      enableColumnFilter: true
    }

    column value #guest_name {
      label: "guest name"
      value: :guest_name
      enableColumnFilter: true
    }

    column value #CustomerPhoneNumber {
      label: "Customer Phone Number"
      value: :CustomerPhoneNumber
      enableColumnFilter: true
    }
    column value #TourSubTotal {
      label: "Tour Sub Total"
      value: :TourSubTotal
      enableColumnFilter: true
    }

    navigateTo: page_Indiv_Survey_Response
  } //end widget
} // end page
page #page_KSCVCResponses {

  label: "Kennedy Space Center - Response Details"

  hide: false
  modal: true

  widget table #tableWidget {
    label: "Kennedy Space Center Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start

    filter expression #expressionFilter {
      value: surveyDataset:filterMeasure_KSCVCSurvey()
      label: "KSCVC survey Only"
    }

    filter expression {
      value: surveyDataset:filterMeasure_NPSanswered()
      label: "NPS has a value"
    }

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      format: valueDefaultFormatter
      enableColumnFilter: true
    }

    column value #LocationName {
      label: "Location Name"
      value: :LocationName
      enableColumnFilter: true
    }

    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
    }


    column value #SAT {
      label: "Overall Satisfaction"
      value: :SAT
      enableColumnFilter: true
    }

    column value #Value {
      label: "Value"
      value: :Value
      enableColumnFilter: true
    }


    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
    }

    column value #EXPERIENCES {
      label: "EXPERIENCES"
      value: :EXPERIENCES
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_attractions {
      label: "Sat-Attractions"
      value: :SAT_EXPERIENCES.attractions
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_bus {
      label: "Sat-Bus Tour"
      value: :SAT_EXPERIENCES.bus
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_premiums {
      label: "Sat-Premiums"
      value: :SAT_EXPERIENCES.premiums
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_restaurants {
      label: "Sat-Restaurants"
      value: :SAT_EXPERIENCES.restaurants
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_shops {
      label: "Sat-Shops"
      value: :SAT_EXPERIENCES.shops
      enableColumnFilter: true
    }

    column value #SAT_EXPERIENCES_rides {
      label: "Sat-Rides"
      value: :SAT_EXPERIENCES.rides
      enableColumnFilter: true
    }


    column value #ATTRACTIONS_SEEN {
      label: "ATTRACTIONS SEEN"
      value: :ATTRACTIONS_SEEN
      enableColumnFilter: true
    }


    column value #ATTRACT_INSERT {
      label: "ATTRACTION INSERT"
      value: :ATTRACT_INSERT
      enableColumnFilter: true
    }

    column value #DRILL_ATTRACTION_cleanliness {
      label: "Sat-Attraction Cleanliness"
      value: :DRILL_ATTRACTION.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_ATTRACTION_quality {
      label: "Sat-Attraction Quality"
      value: :DRILL_ATTRACTION.quality
      enableColumnFilter: true
    }
    column value #DRILL_ATTRACTION_staff {
      label: "Sat-Attraction Staff"
      value: :DRILL_ATTRACTION.staff
      enableColumnFilter: true
    }
    column value #DRILL_BUS_cleanarea {
      label: "Sat-Bus Tours-Waiting Area"
      value: :DRILL_BUS.cleanarea
      enableColumnFilter: true
    }
    column value #DRILL_BUS_cleanbus {
      label: "Sat-Bus Tours-Clean"
      value: :DRILL_BUS.cleanbus
      enableColumnFilter: true
    }
    column value #DRILL_BUS_quality {
      label: "Sat-Bus Tours-Quality"
      value: :DRILL_BUS.quality
      enableColumnFilter: true
    }
    column value #DRILL_BUS_staff {
      label: "Sat-Bus Tours-Staff"
      value: :DRILL_BUS.staff
      enableColumnFilter: true
    }
    column value #DRILL_BUS_waitime {
      label: "Sat-Bus Tours-Wait Time"
      value: :DRILL_BUS.waitime
      enableColumnFilter: true
    }

    column value #RESTAURANT_INSERT {
      label: "RESTAURANT_INSERT"
      value: :RESTAURANT_INSERT
      enableColumnFilter: true
    }

    column value #DRILL_RESTAURANT_cleanliness {
      label: "Restaurant-Cleanliness"
      value: :DRILL_RESTAURANT.cleanliness
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_kiosk {
      label: "Restaurant-Kiosk"
      value: :DRILL_RESTAURANT.kiosk
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_quality {
      label: "Restaurant-Quality of food/bev"
      value: :DRILL_RESTAURANT.quality
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_speed {
      label: "Restaurant-Speed of service"
      value: :DRILL_RESTAURANT.speed
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_staff {
      label: "Restaurant-Staff"
      value: :DRILL_RESTAURANT.staff
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_value {
      label: "Restaurant-Value"
      value: :DRILL_RESTAURANT.value
      enableColumnFilter: true
    }
    column value #DRILL_RESTAURANT_variety {
      label: "Restaurant-Variety"
      value: :DRILL_RESTAURANT.variety
      enableColumnFilter: true
    }

    column value #RESTAURANT_COMMENTS {
      label: "RESTAURANT_COMMENTS"
      value: :RESTAURANT_COMMENTS
      enableColumnFilter: true
    }

    column value #PREMIUM_PURCHASED {
      label: "PREMIUM_PURCHASED"
      value: :PREMIUM_PURCHASED
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_foodquality {
      label: "Sat-Premium-Food Quality"
      value: :DRILL_PREMIUM.foodquality
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_quality {
      label: "Sat-Premium-Tour Quality"
      value: :DRILL_PREMIUM.quality
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_staff {
      label: "Sat-Premium-Staff"
      value: :DRILL_PREMIUM.staff
      enableColumnFilter: true
    }
    column value #DRILL_PREMIUM_value {
      label: "Sat-Premium-Value"
      value: :DRILL_PREMIUM.value
      enableColumnFilter: true
    }
    column value #SHOPS_VISITED {
      label: "SHOPS_VISITED"
      value: :SHOPS_VISITED
      enableColumnFilter: true
    }
    column value #SHOPS_INSERT {
      label: "SHOPS_INSERT"
      value: :SHOPS_INSERT
      enableColumnFilter: true
    }
    column value #PURCHASE {
      label: "Purchase Made"
      value: :PURCHASE
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_shopsat {
      label: "Sat-Shops-OSAT"
      value: :DRILL_SHOPS.shopsat
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_merch {
      label: "Sat-Shops-Merch Quality"
      value: :DRILL_SHOPS.merch
      enableColumnFilter: true
    }

    column value #DRILL_SHOPS_speed {
      label: "Sat-Shops-Speed of Checkout"
      value: :DRILL_SHOPS.speed
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_staff {
      label: "Sat-Shops-Staff"
      value: :DRILL_SHOPS.staff
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_value {
      label: "Sat-Shops-Value"
      value: :DRILL_SHOPS.value
      enableColumnFilter: true
    }
    column value #DRILL_SHOPS_variety {
      label: "Sat-Shops-Variety"
      value: :DRILL_SHOPS.variety
      enableColumnFilter: true
    }

    column value #Problem {
      label: "Problem"
      value: :PROBLEM
      enableColumnFilter: true
    }
    column value #PROB_REPORTED {
      label: "Problem Reported"
      value: :PROB_REPORTED
      enableColumnFilter: true
    }
    column value #RESOLUTION_SAT {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    column value #CONTACT_REQUESTED {
      label: "Contact Requested"
      value: :CONTACT
      enableColumnFilter: true
    }
    column value #CONTACT_PREF {
      label: "Method of Contact"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_name {
      label: "Contact Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_phone {
      label: "Contact Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_email {
      label: "Contact Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #PROBLEM_DETAIL {
      label: "Problem Detail"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #TEAM_REC {
      label: "Team Recognition"
      value: :TEAM_REC
      enableColumnFilter: true
    }
    column value #TEAM_MEMBER {
      label: "Team Member"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #RECOG_DETAIL {
      label: "Team Recognition Detail"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }
    //start demos
    column value #REGION {
      label: "REGION"
      value: :REGION
      enableColumnFilter: true
    }
    column value #GENDER {
      label: "GENDER"
      value: :GENDER
      enableColumnFilter: true
    }
    column value #AGE {
      label: "AGE"
      value: :AGE
      enableColumnFilter: true
    }
    column value #INCOME {
      label: "INCOME"
      value: :INCOME
      enableColumnFilter: true
    }
    column value #UNDER_18_KIDS {
      label: "UNDER_18_KIDS"
      value: :UNDER_18_KIDS
      enableColumnFilter: true
    }
    column value #EDUCATION {
      label: "EDUCATION"
      value: :EDUCATION
      enableColumnFilter: true
    }
    column value #ETHNICITY {
      label: "ETHNICITY"
      value: :ETHNICITY
      enableColumnFilter: true
    }
    column value #NO_VISITS {
      label: "NO_VISITS"
      value: :NO_VISITS
      enableColumnFilter: true
    }
    column value #AWARENESS {
      label: "AWARENESS"
      value: :AWARENESS
      enableColumnFilter: true
    }
    column value #KSC_COMPANIONS {
      label: "KSC_COMPANIONS"
      value: :KSC_COMPANIONS
      enableColumnFilter: true
    }
    column value #TOTAL_PARTY {
      label: "TOTAL_PARTY"
      value: :TOTAL_PARTY
      enableColumnFilter: true
    }

    column value #ACCOMMODATIONS {
      label: "ACCOMMODATIONS"
      value: :ACCOMMODATIONS
      enableColumnFilter: true
    }
    column value #KSC_LOCATION {
      label: "LOCATION"
      value: :LOCATION
      enableColumnFilter: true
    }
    column value #OTHER_ATTRACTIONS {
      label: "OTHER_ATTRACTIONS"
      value: :OTHER_ATTRACTIONS
      enableColumnFilter: true
    }
    column value #NO_VACATIONS {
      label: "NO_VACATIONS"
      value: :NO_VACATIONS
      enableColumnFilter: true
    }

  //start BG info
    column value #email {
      label: "email"
      value: :email
      enableColumnFilter: true
    }

    column value #Postal {
      label: "Postal"
      value: :Postal
      enableColumnFilter: true
    }

    column value #guest_name {
      label: "guest_name"
      value: :guest_name
      enableColumnFilter: true
    }
    column value #TransactionID {
      label: "TransactionID"
      value: :TransactionID
      enableColumnFilter: true
    }

    column date #YieldDateTime {
      label: "YieldDateTime"
      value: :YieldDateTime
      enableColumnFilter: true
    }
    column value #CountryName {
      label: "CountryName"
      value: :CountryName
      enableColumnFilter: true
    }
    column value #CompanyID {
      label: "CompanyID"
      value: :CompanyID
      enableColumnFilter: true
    }
    column value #NodeNo {
      label: "NodeNo"
      value: :NodeNo
      enableColumnFilter: true
    }
    column value #SellingPrice {
      label: "SellingPrice"
      value: :SellingPrice
      enableColumnFilter: true
    }
    column value #UseNo {
      label: "UseNo"
      value: :UseNo
      enableColumnFilter: true
    }

    navigateTo: page_Indiv_Survey_Response
  } //end widget
} // end page
page #page_DNListensResponses {

  label: "DN Listens - Response Details"
  hide: false
  modal: true

  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_DNListensSurvey()
    label: "DN Listens Only"
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  widget table #tableWidget {
    label: "Travel Hospitality - Responses"
    size: "large"
    table: :
    paginationType: paging
    sortOrder: descending
    sortColumn: interview_start
    rowsPerPage: 100, 500, 1000

    column date #interview_start {
      label: "Interview Date"
      value: :interview_start
      enableColumnFilter: true
    }
    column value #interview_status {
      label: "Interview Status"
      value: :status
      enableColumnFilter: true
    }
    column value #SurveyType {
      label: "Survey Type (DN Listens)"
      value: :SurveyType
      enableColumnFilter: true
    }
    column value #LocationName {
      label: "Location Name"
      //value: :LocationFinal
      value: demote(SitesHierarchy:language_text, surveyDataset:)
      enableColumnFilter: true
    }
    column date #VISIT_DATE {
      label: "Visit Date"
      value: :VISIT_DATE
      enableColumnFilter: true
    }
    column value #TIME_OF_VISIT {
      label: "Time of Visit"
      value: :TIME_OF_VISIT
      enableColumnFilter: true
    }
    column value #STORE_INFO {
      label: "Store Info"
      value: :STORE_INFO
      enableColumnFilter: true
    }

    column value #StateProvince {
      label: "State / Province"
      value: :StateProvince
      enableColumnFilter: true
    }
    column value #NPS {
      label: "NPS"
      value: :NPS
      enableColumnFilter: true
    }

    column value #SAT {
      label: "Overall Satisfaction"
      value: :SAT
      enableColumnFilter: true
    }

    column value #SAT_DRIVERS_quality {
      label: "Food quality"
      value: :SAT_DRIVERS.quality
      enableColumnFilter: true
    }

    column value #SAT_DRIVERS_speed {
      label: "Speed of service"
      value: :SAT_DRIVERS.speed
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_staff {
      label: "Staff"
      value: :SAT_DRIVERS.staff
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_value {
      label: "Value"
      value: :SAT_DRIVERS.value
      enableColumnFilter: true
    }
    column value #SAT_DRIVERS_variety {
      label: "Variety of items available"
      value: :SAT_DRIVERS.variety
      enableColumnFilter: true
    }

    column value #VISIT_COMMENTS {
      label: "Visit Comments"
      value: :VISIT_COMMENTS
      enableColumnFilter: true
    }

    column value #Problem {
      label: "Problem"
      value: :PROBLEM
      enableColumnFilter: true
    }
    column value #PROB_REPORTED {
      label: "Problem Reported"
      value: :PROB_REPORTED
      enableColumnFilter: true
    }
    column value #RESOLUTION_SAT {
      label: "Problem Resolution Sat"
      value: :RESOLUTION_SAT
      enableColumnFilter: true
    }
    column value #CONTACT_REQUESTED {
      label: "Contact Requested"
      value: :CONTACT
      enableColumnFilter: true
    }
    column value #CONTACT_PREF {
      label: "Method of Contact"
      value: :CONTACT_PREF
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_name {
      label: "Contact Name"
      value: :CONTACT_INFO.name
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_phone {
      label: "Contact Phone"
      value: :CONTACT_INFO.phone
      enableColumnFilter: true
    }
    column value #CONTACT_INFO_email {
      label: "Contact Email"
      value: :CONTACT_INFO.email
      enableColumnFilter: true
    }
    column value #PROBLEM_DETAIL {
      label: "Problem Detail"
      value: :PROBLEM_DETAIL
      enableColumnFilter: true
    }
    column value #TEAM_REC {
      label: "Team Recognition"
      value: :TEAM_REC
      enableColumnFilter: true
    }
    column value #TEAM_MEMBER {
      label: "Team Member"
      value: :TEAM_MEMBER
      enableColumnFilter: true
    }
    column value #RECOG_DETAIL {
      label: "Team Recognition Detail"
      value: :RECOG_DETAIL
      enableColumnFilter: true
    }

    column value #LOI {
      label: "LOI"
      value: :LOI
      enableColumnFilter: true
    }

    navigateTo: page_Indiv_Survey_Response
  } //end widget
} // end page
page #page_ResponseDiagnostics {

  label: "Response Diagnostics"
  widget headline #headlineWidget {
    size: large

    tile markdown #markdownTile_2 {
      value: "# Response Diagnostics

***Note: DN Listens survey results are not included on this page.***"

    } //end widget
    label: "Voice of Guest Dashboard"
  }

//  hide: true
  modal: false
  ignoreFilters: reportingPeriodFilter, f_Surveys, f_Location
  overrideFilter date {
    dateVariables: @reportConfig.InvitedDate
  }

  access rules {
    rule claim {
      name: "UserLevel"
      value: "Power User"
    }
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  layoutArea toolbar {
    useDynamicFilters: true
    filter date {
      dateVariables: @reportConfig.InvitedDate
      dateOption YearToDate {
        label: "Year to date"
        selected: true
      }
      label: "Invited Date"
    }

    filter multiselect #f_SurveysRespData {
      optionsFrom: surveyDataset.respondent:survey_pid
      label: "Survey Name"
    }

    filter multiselect #f_LocationResp {
      optionsFrom: surveyDataset.respondent:LocationName
      label: "Location"
    }

  } //end widget
  widget kpi #kpiWidget_RespRate {
    label: "Overall Response Rate"
   // label: "Response Rate (Does not work with filters applied) "
   // hide: true
    filter expression {
      value: _not(IN(:survey_pid, @reportConfig.surveypid_dnlistens))
  //not dn listens

    }
    tile kpi #kpiTile {

      value: count(@reportConfig.nps_qid) / count(.respondent:, @reportConfig.emailsSent) * 100

      format: oneDecimalPercent
      min: 0
      max: 100
      //target: 25
      showRange: true
      navigateTo: page_KPIBreakdowns
    }

    tile value {
      label: "No. Invited"
      value: count(.respondent:, @reportConfig.emailsSent)
      format: noDecimalNumber
    }

    tile value {
      label: "No. Responses"
      value: count(@reportConfig.nps_qid)
      format: noDecimalNumber

    }

    infobox {
      label: "Response Rate"
      info: @reportConfig.ResponseRateNote
    }
    description: "This widget does not include DN Listens survey which is an open survey"
  } // end widget
  widget chart #chartWidget_RespRateTrends {
    label: "Response Rate Trends"
    size: medium
    legend: "none"
    palette: survey_metrics_palette
    removeEmptyCategories: true
    removeEmptySeries: true
    ignoreFilters: reportingPeriodFilter
   //   significanceTesting: true    
   // hide: true
    filter expression {
      value: @Timeframe_Selector_RR.selected.selectFilter
    }

    filter expression {
      value: _not(IN(:survey_pid, @reportConfig.surveypid_dnlistens))
  //not dn listens

    }
 //here is an inline selector
    select #Timeframe_Selector_RR {
      label: "Select a Timeframe"

      options: @valueSet_date_ranges_RR.items

    } // end selector
    series {
      value: count(@reportConfig.nps_qid) / count(.respondent:, @reportConfig.emailsSent) * 100
        //    value: count(@reportConfig.nps_qid)

      format: oneDecimalPercent
     // format: twoDecimalNumber   
      label: "Response Rate"
      chart bar #undefined {
        maxBarSize: 100

      }
      //percentOver: "series"
    }

    category date #cutByDate {
      value: @reportConfig.InvitedDate
      breakdownBy: @Timeframe_Selector_RR.selected.selectBreakdownBy
      label: "Invited date"
      //format: dateDefaultFormatter
    }

    axis category #categoryAxis {
      orientation: "-45"
      interval: "all"
      label: "Invited date"
      textSize: 80
    }
    axis primary #primaryAxis {
      minValue: 0
      format: noDecimalPercent
      label: "Response Rate (%)"
    }

    axis secondary {
    }

    infobox {
      label: "Response Rate"
      info: "NOTE: Response Rate = (# Respondents who answered the first question) / (# Invited)"
    }
    base #base {
      value: count(.respondent:, @reportConfig.emailsSent)
      format: baseNumberFormatter
    }


    description: "This widget does not include DN Listens survey which is an open survey"
  } // end widget
  widget dataGrid #dataGridWidget_2 {
    label: "Response Rates by Location"
    size: halfwidth
    ignoreFilters: f_Location, reportingPeriodFilter
    removeEmptyRows: true
    showLegend: false


    filter expression {
      value: _not(IN(:survey_pid, @reportConfig.surveypid_dnlistens))
  //not dn listens

    }
 //here is an inline selector
    select #Timeframe_Selector_RR {
      label: "Select a Timeframe"

      options: @valueSet_date_ranges_RR.items

    } // end selector
    row comparison {
      reportingHierarchy: LocationsBySurveyHierarchy

    }

    column {

      cell {
        value: count(@reportConfig.nps_qid) / count(.respondent:, @reportConfig.emailsSent) * 100
        format: oneDecimalPercent
        extraValue: count(.respondent:, @reportConfig.emailsSent)
        extraValueFormat: noDecimalNumber
      }

      label: "Response Rate"
    }
    column {
      label: "Response Rate Trends"

      cell microchart {

        value: count(@reportConfig.nps_qid) / count(.respondent:, @reportConfig.emailsSent) * 100

        format: oneDecimalPercent
        useOnlyExistingColumns: true
        extraValue: count(.respondent:, @reportConfig.emailsSent)
        extraValueFormat: noDecimalNumber
        breakdownBy date {
          value: @reportConfig.InvitedDate
          breakdownBy: @Timeframe_Selector_RR.selected.selectBreakdownBy

         // format: dateFormatDay
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

  } // end widget
  widget chart #chartWidget_6 {
    label: "Response Rate By Survey"
    size: medium
    legend: "none"
    palette: survey_metrics_palette
    removeEmptyCategories: true
    removeEmptySeries: true
    ignoreFilters: reportingPeriodFilter
   //   significanceTesting: true    


    filter expression {
      value: _not(IN(:survey_pid, @reportConfig.surveypid_dnlistens))
  //not dn listens

    }

    series {
      value: count(@reportConfig.nps_qid) / count(.respondent:, @reportConfig.emailsSent) * 100
        //    value: count(@reportConfig.nps_qid)

      format: oneDecimalPercent
     // format: twoDecimalNumber   
      label: "Response Rate"
      chart bar #undefined {
        maxBarSize: 75

      }
      //percentOver: "series"
    }

    category cut {
      value: .respondent:survey_pid

    }

    axis category #categoryAxis {
      orientation: "0"
      interval: "all"
      label: "Survey Name"
      textSize: 55
    }
    axis primary #primaryAxis {
      minValue: 0
      format: noDecimalPercent
      label: "Response Rate (%)"
    }

    axis secondary {
      hide: true
    }

    infobox {
      label: "Response Rate"
      info: "NOTE: Response Rate = (# Respondents who answered the first question) / (# Invited)"
    }
    base #base {
      value: count(.respondent:, @reportConfig.emailsSent)
      format: baseNumberFormatter
    }

    description: "This widget does not include DN Listens survey which is an open survey"
  } // end widget
  widget chart #chartWidget {
    label: "Responses By Survey"
    //animation: true
    size: medium
    //gridLines: both
    legend: bottomCenter
    palette: survey_metrics_palette
    removeEmptyCategories: true
    removeEmptySeries: true

    filter expression {
      value: IN(.respondent:responseStatus, "c", "i")

    }
    series {
      value: count(.respondent:responseStatus)
      format: noDecimalNumber
      breakdownBy cut {
        value: .respondent:responseStatus
      }
      chart bar {
        mode: stacked
        maxBarSize: 75
      }
    }
    axis secondary {
      //minValue: 0
     // maxValue: 100
    }

    category cut {
      value: :survey_pid

    }
    //ignoreFilters: period
    axis category #categoryAxis {
      label: "Survey Name"
      textSize: 55
    }
    axis primary #primaryAxis {
      format: noDecimalNumber
    }
    //navigateTo: group_drilldown
    base #base {
      value: count(.respondent:responseStatus)
      format: baseNumberFormatter
    }
  } // end widget
  widget dataGrid #dataGridWidget_5 {
    label: "Daily Response Status (Last 7 days)"
    size: large
    ignoreFilters: f_Location, reportingPeriodFilter
    removeEmptyRows: true
    showLegend: false
    filter expression {
      value: InDay(surveyDataset.respondent:CreatedDate, -6, 0)
    }

    view comparativeStatistic #zerosView {
      valueColorFormatter: text_zeros_formatter
      backgroundColorFormatter: background_zeros_formatter
    }

    row comparison {
      reportingHierarchy: LocationsBySurveyHierarchy
    }

    column {
      label: "Num Loaded Last 7 days"

      cell microchart {

        value: count(surveyDataset.respondent:CreatedDate)
        format: noDecimalNumber
        useOnlyExistingColumns: true

        breakdownBy date {
          value: surveyDataset.respondent:CreatedDate
          breakdownBy: calendarDate
          format: dateFormatDay
        }

        microchart line {
          showDots: true
          showTooltip: true
          color: #1D78BA
        }
      }

    }

    column cutByDate {
      value: surveyDataset.respondent:CreatedDate
      breakdownBy: calendarDate
      format: dateFormatDay
    //  movingAverageStart: "7 days"
      sortOrder: descending
      total: none
      column {

        cell {
          value: count(surveyDataset.respondent:CreatedDate)
          format: noDecimalNumber
          view: zerosView
          navigateTo: page_RespondentDetails
        }
        label: "Num Loaded"
      }
      column cut {
        value: surveyDataset.respondent:responseStatus
        total: none
        categories: "'c','i'"
        cell {
          value: count(surveyDataset.respondent:responseStatus)
          format: noDecimalNumber

        }
      }
    }

    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: copy_of_sentimentindicatortext
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }
  } // end widget
  widget chart #chartWidget_2 {
    label: "Daily Responses (Last 45 days)"
    //animation: true
    size: large
    //gridLines: both
    legend: bottomCenter
    palette: survey_metrics_palette
    removeEmptyCategories: true
    removeEmptySeries: true
    //experimentalTooltip: true
    chartMargin {
      bottom: 10
    }
    filter expression {
      value: InDay(@reportConfig.intvdate, -44, 0)

    }
    filter expression {
      value: IN(.respondent:responseStatus, "c", "i")

    }

    series {
      value: count(.respondent:responseStatus)
      format: noDecimalNumber

      breakdownBy cut {
        value: .respondent:responseStatus
      }
      chart bar {
        mode: stacked
      }
    }
    axis secondary {
     // minValue: 0
     // maxValue: 100
    }

    category date {

      value: @reportConfig.intvdate
      //breakdownBy: calendarMonth
      breakdownBy: calendarDate
      label: "Date"
      format: dateFormatDay
    }

    axis category #categoryAxis {
      orientation: "-45"
      label: "Interview Date"
    }
    axis primary #primaryAxis {
      format: noDecimalNumber
    }

  }
  widget chart #chartWidget_3 {
    label: "By Device Type"
    layout: "horizontal"
    legend: bottomCenter
    size: small
    palette: survey_metrics_palette

    removeEmptyCategories: true

    chart bar {
      mode: clustered
    }

    series {
      value: count(surveyDataset:)
      percentOver: series
      format: oneDecimalPercent
      chart bar #barChart {
        mode: "clustered"
        maxBarSize: 50
      }
      breakdownBy cut #cutBreakdownby {
        value: surveyDataset:lastdevicetype
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    removeEmptySeries: true


    base #base {
      value: count(surveyDataset:lastdevicetype)
      format: baseNumberFormatter
    }

  } // end widget
  widget chart #chartWidget_LOI {
    label: "Length of Interview By Survey (median)"

    size: medium

    legend: "none"
    palette: survey_metrics_palette
    removeEmptyCategories: true
    removeEmptySeries: true


    series {
      label: "Median LOI (in mins)"
      value: median(:LOI)
      format: twoDecimalNumber
      chart bar {

        maxBarSize: 65
      }
    }
    axis secondary {
      //minValue: 0
     // maxValue: 100
    }

    category cut {
      value: :survey_pid

    }

    axis category #categoryAxis {

      label: "Survey Name"
    }
    axis primary #primaryAxis {
      format: noDecimalNumber
      label: "LOI (in minutes)"
      minValue: 0
    }

    base #base {
      value: count(:survey_pid)
      format: baseNumberFormatter
    }
  } // end widget
  config layout #layoutConfig {
    horizontalAlignmentMode: "fourColumnsCentered"
  }
} // end page
page #page_Demos {
  label: "Demographics"
  widget markdown #markdownWidget {
    markdown: "# **Survey Demographics**
### This page provides a breakdown of key guest demographic categories; this can be helpful in understanding who is responding to our surveys.

"
    size: large
  }

  widget chart #chartWidget_Demos_Region {
    label: "Region"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

//hide: IIF(count(surveyDataset:status = "complete") < 1, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :REGION
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Region_Alt {
    label: "Region (Australia locations)"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

//hide: IIF(count(surveyDataset:status = "complete") < 1, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :REGION_ALPHA
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Gender {
    label: "Gender"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :GENDER
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Age {
    label: "Age"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :AGE
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Income {
    label: "Income"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :INCOME
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_NumKids {
    label: "No. of Kids Under 18"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :UNDER_18_KIDS
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Education {
    label: "Education"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :EDUCATION
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Ethnicity {
    label: "Ethnicity"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :ETHNICITY
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_NumVisits {
    label: "Number of Visits"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :NO_VISITS
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Companions {
    label: "Companions on Trip"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :COMPANIONS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #chartWidget_Demos_Leisure {
    label: "Ave No. of Leisure Trips/Yr"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :NO_VACATIONS
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #copy_of_copy_of_chartWidget_Demos_Leisure {
    label: "Survey Source Data (Used for Checking)"
    // suppressRule {
    //   criteria: @reportConfig.suppressCriteriaMin
    // }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 60
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
      minValue: 0
      maxValue: 100
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :combined_sourceid
    }
    chartMargin {
      left: 20
    }
  } // end widget
  modal: true
  hide: false
} // end page
page #page_Demos_Gaming {
  label: "Demographics - Gaming"
  widget markdown #markdownWidget {
    markdown: "# **Survey Demographics**
### This page provides a breakdown of key guest demographic categories; this can be helpful in understanding who is responding to our surveys.

"
    size: large
  }

  widget chart #chartWidget_Demos_Region {
    label: "Region"
    // suppressRule {
    //   criteria: @reportConfig.suppressCriteriaMin
    // }
//hide: count(surveyDataset:status = "complete") > 1
//hide: IIF(count(surveyDataset:status = "complete") < 1, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :REGION
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Gender {
    label: "Gender"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :GENDER
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Age {
    label: "Age"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :AGE
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Income {
    label: "Income"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :INCOME
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_NumKids {
    label: "No. of Kids Under 18"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :UNDER_18_KIDS
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Education {
    label: "Education"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :EDUCATION
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Ethnicity {
    label: "Ethnicity"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :ETHNICITY
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Ethnicity_AUS {
    label: "Ethnicity (Australia locations)"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :ETHNICITY_AUS
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Companions {
    label: "Companions on Trip"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :COMPANIONS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #copy_of_chartWidget_Demos_Companions {
    label: "Total People In Party"
    // suppressRule {
    //   criteria: @reportConfig.suppressCriteriaMin
    // }
    //hide:@reportConfig.suppressCriteriaMin
    //hide: IIF(count(:) = 0, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :TOTAL_PARTY
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #copy_of_copy_of_chartWidget_Demos_Companions {
    label: "Time of Gaming Visit"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :TIME_OF_GAMING_VISIT
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #copy_of_chartWidget_Demos_Leisure_2 {
    label: "Did You Win or Lose on This Trip?"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :WIN_LOSE
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #copy_of_copy_of_chartWidget_Demos_Leisure_2 {
    label: "Did Visit Include a Special Event?"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :SPEC_EVENT
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget comments #copy_of_copy_of_commentsWidget {
    label: "Other Special Event"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Other Type of Special Event"
      filter expression #excludeBlankResponses {
        value: :SPEC_EVENT.98$other != ""
      }
      comment: :SPEC_EVENT.98$other
    }
    size: "medium"
    table: :
    column value #valueColumn {
      label: "Gaming Facility"
      value: :casino_name
    }
  }
  widget chart #copy_of_copy_of_copy_of_chartWidget_Demos_Leisure_2 {
    label: "Comps Received During Visit"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :COMPS
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget comments #copy_of_commentsWidget {
    label: "Other Types of Comps Received"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Other Redemption Type"
      filter expression #excludeBlankResponses {
        value: :COMPS.98$other != ""
      }
      comment: :COMPS.98$other
    }
    size: "medium"
    table: :
    column value #valueColumn {
      label: "Gaming Facility"
      value: :casino_name
    }
  }
  widget chart #copy_of_copy_of_copy_of_copy_of_chartWidget_Demos_Leisure_2 {
    label: "Points Redeemed For..."
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :REDEMPTION
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget comments #commentsWidget {
    label: "Other Redemption Used"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Other Redemption Type"
      filter expression #excludeBlankResponses {
        value: :REDEMPTION.98$other != ""
      }
      comment: :REDEMPTION.98$other
    }
    size: "medium"
    table: :
    column value #valueColumn {
      label: "Gaming Facility"
      value: :casino_name
    }
  }
  widget chart #copy_of_copy_of_chartWidget_Demos_Leisure {
    label: "Survey Source Data (Used for Checking)"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: large
    layout: "vertical"
    category cut #cutCategory {
      value: :combined_sourceid
    }
    chartMargin {
      left: 20
    }
  } // end widget
  modal: true
  hide: false
} // end page
page #page_Demos_KSCVC {
  label: "Demographics - Kennedy Space Center"

  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_KSCVCSurvey()
    label: "KSCVC survey Only"
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  widget markdown #markdownWidget {
    markdown: "# **Survey Demographics - Kennedy Space Center**
### This page provides a breakdown of key guest demographic categories; this can be helpful in understanding who is responding to our surveys.

"
    size: large
  }

  widget chart #chartWidget_Demos_Region {
    label: "Region"
    // suppressRule {
    //   criteria: @reportConfig.suppressCriteriaMin
    // }
//hide: count(surveyDataset:status = "complete") > 1
//hide: IIF(count(surveyDataset:status = "complete") < 1, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :REGION
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Gender {
    label: "Gender"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :GENDER
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Age {
    label: "Age"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :AGE
      //sortOrder: descending
      //sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Income {
    label: "Income"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :INCOME
      //sortOrder: descending
      //sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_NumKids {
    label: "No. of Kids Under 18"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :UNDER_18_KIDS
      //sortOrder: descending
      //sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Education {
    label: "Education"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :EDUCATION
      //sortOrder: descending
      //sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Ethnicity {
    label: "Ethnicity"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :ETHNICITY
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Awareness {
    label: "Methods of Awareness"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :AWARENESS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #chartWidget_Demos_ksc_companions {
    label: "Travel Companions - This Trip"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :KSC_COMPANIONS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #chartWidget_Demos_NumInParty {
    label: "Total People In Party"
    // suppressRule {
    //   criteria: @reportConfig.suppressCriteriaMin
    // }
    //hide:@reportConfig.suppressCriteriaMin
    //hide: IIF(count(:) = 0, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :TOTAL_PARTY
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #chartWidget_Demos_NumVisits {
    label: "No. of Visits"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :NO_VISITS
     // sortOrder: descending
      //sortBy: "series"
    }
    chartMargin {
      left: 40
    }
  } // end widget
  widget chart #chartWidget_Demos_FlaAccommodations {
    label: "Florida Accommodations"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :ACCOMMODATIONS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_FlaLocation {
    label: "Florida Location"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :LOCATION
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_OtherAttractions {
    label: "Other Attractions Visited"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cutByMulti #cutCategory {
      value: :OTHER_ATTRACTIONS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_NumVacations {
    label: "Typical No. of Trips/Yr"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :NO_VACATIONS
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Survey {
    label: "Survey Source Data (Used for Checking)"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: large
    layout: "vertical"
    category cut #cutCategory {
      value: :survey_name
    }
    chartMargin {
      left: 20
    }
  } // end widget
  modal: true
  hide: false
} // end page
page #page_Demos_LizardIsland {
  label: "Demographics - Lizard Island"

  filter expression #expressionFilter {
    value: surveyDataset:filterMeasure_LizardIslandSurvey()
    label: "Lizard Island survey only"
  }

  filter expression {
    value: surveyDataset:filterMeasure_NPSanswered()
    label: "NPS has a value"
  }

  widget markdown #markdownWidget {
    markdown: "# **Survey Demographics - Lizard Island**
### This page provides a breakdown of key guest demographic categories; this can be helpful in understanding who is responding to our surveys.

"
    size: large
  }

  widget chart #chartWidget_Demos_Region {
    label: "Region"
    // suppressRule {
    //   criteria: @reportConfig.suppressCriteriaMin
    // }
//hide: count(surveyDataset:status = "complete") > 1
//hide: IIF(count(surveyDataset:status = "complete") < 1, true, false)
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :REGION_ALPHA
      sortOrder: descending
      sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Age {
    label: "Age"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }

    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
        maxBarSize: 65
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: halfwidth
    layout: "horizontal"
    category cut #cutCategory {
      value: :AGE
      //sortOrder: descending
      //sortBy: "series"
    }
    chartMargin {
      left: 20
    }
  } // end widget
  widget chart #chartWidget_Demos_Survey {
    label: "Survey Source Data (Used for Checking)"
    suppressRule {
      criteria: @reportConfig.suppressCriteriaMin
    }
    series #series {
      chart bar #barChart {
        showBase: true
        showValue: true
      }
      value: count(:)
      percentOver: "categories"
      format: oneDecimalPercent
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      label: "Percentage"
      format: noDecimalPercent
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: large
    layout: "vertical"
    category cut #cutCategory {
      value: :survey_name
    }
    chartMargin {
      left: 20
    }
  } // end widget
  modal: true
  hide: false
} // end page
page #page_RespondentDetails {
  label: "Respondent Details"
  widget table #tableWidget {
    label: "Respondent Table"
    size: "large"
    table: .respondent:
    column date #CreatedDate {
      label: "CreatedDate"
      value: .respondent:CreatedDate
      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "survey_rid"
      value: .respondent:survey_rid
      enableColumnFilter: true
    }
    column value #valueColumn_3 {
      label: "survey_name"
      value: .respondent:survey_name
      enableColumnFilter: true
    }
    column value #valueColumn_4 {
      label: "survey_pid"
      value: .respondent:survey_pid
      enableColumnFilter: true
    }
    column value #valueColumn_5 {
      label: "combined_sourceid"
      value: .respondent:combined_sourceid
      enableColumnFilter: true
    }
    column value #valueColumn_6 {
      label: "combined_sourceid_text"
      value: .respondent:combined_sourceid_text
      enableColumnFilter: true
    }
    sortColumn: CreatedDate
    sortOrder: descending
  } //end widget
  hide: false
  modal: true
} //end page
page #dd_SentimentComments_Lodging {
  modal: true
  hide: false
  label: "Comments Drilldown - Lodging"
  modalSize: large

  widget comments #comments_Lodging {

    table: textAnalyticsDataset_Lodging.overallScore:
    label: "Comments Drilldown - Lodging"
    size: large
    showHeader: true
    sortOrder: descending
    sortColumn: comments
    headerNumberOfLines: 3

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response_TA

    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
      fontSize: medium
    }

    group question {
      label: "All Comments"
      comment: textAnalyticsDataset_Lodging.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Lodging.overallScore:text != ""
      }
    }
    column response #comments {
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta
      view: viewComments
      enableColumnFilter: true
    }
    column value #valueColumn_OpenEnds {
      label: "Comment Field"
      value: textAnalyticsDataset_Lodging.overallScore:variable
      enableColumnFilter: true
      width: 125px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }


    column metric #metricColumn_overall_sentiment {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Lodging:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Lodging:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 150px
    }


    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    // column metric #metricColumn_NPS {
    //   label: "NPS"
    //   value: score(@reportConfig.nps_qid_ta)
    //   enableColumnFilter: true
    //   //filterable: true
    //   width: 125px
    //   align: center
    //   view: colorcoding


    // }

    // column metric #metricColumn_OSAT {
    //   label: "SAT"
    //   value: score(@reportConfig.osat_qid_ta)
    //   enableColumnFilter: true
    //   width: 125px
    //   align: center
    //   view: colorcoding_5pt
    // }

    // column metric #metricColumn_Value {
    //   label: "Value"
    //   value: score(@reportConfig.value_qid_ta)
    //   enableColumnFilter: true
    //   width: 125px
    //   align: center
    //   view: colorcoding_5pt
    // }

    view comment #viewComments {
      lines: 10
    }

  } // end widget
} // end page
page #dd_SentimentComments_Gaming {
  modal: true
  hide: false
  label: "Comments Drilldown - Gaming"
  modalSize: large

  widget comments #comments_Gaming {

    table: textAnalyticsDataset_Gaming.overallScore:
    label: "Comments Drilldown - Gaming"
    size: large
    showHeader: true
    sortOrder: descending
    sortColumn: comments
    headerNumberOfLines: 3

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response_TA

    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
      fontSize: medium
    }

    group question {
      label: "All Comments"
      comment: textAnalyticsDataset_Gaming.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Gaming.overallScore:text != ""
      }
    }
    column response #comments {
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta
      view: viewComments
      enableColumnFilter: true
    }
    column value #valueColumn_OpenEnds {
      label: "Comment Field"
      value: textAnalyticsDataset_Gaming.overallScore:variable
      enableColumnFilter: true
      width: 125px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #LoyaltyTier {
      label: "Loyalty Tier"
      value: surveyDataset:rank_description
      //value: surveyDataset:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 100px
    }

    column metric #metricColumn_overall_sentiment {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Gaming:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Gaming:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 150px
    }


    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    column metric #metricColumn_NPS {
      label: "NPS"
      value: score(@reportConfig.nps_qid_ta)
      enableColumnFilter: true
      //filterable: true
      width: 125px
      align: center
      view: colorcoding
      show: false

    }

    column metric #metricColumn_OSAT {
      label: "SAT"
      value: score(@reportConfig.osat_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false
    }

    column metric #metricColumn_Value {
      label: "Value"
      value: score(@reportConfig.value_qid_ta)
      enableColumnFilter: true
      width: 125px
      align: center
      view: colorcoding_5pt
      show: false

    }

    view comment #viewComments {
      lines: 10
    }

  } // end widget
} // end page
page #dd_SentimentComments_Dining {
  modal: true
  hide: false
  label: "Comments Drilldown - Dining"
  modalSize: large


  widget comments #commentsWidget_Dining {

    table: textAnalyticsDataset_Dining.overallScore:
    label: "Comments Drilldown - Dining"
    size: large
    showHeader: true
    sortOrder: descending
    sortColumn: comments
    headerNumberOfLines: 3

    paginationType: paging
    rowsPerPage: 100, 250, 500, 1000

    navigateTo: page_Indiv_Survey_Response_TA

    view metric #colorcoding {
      backgroundColorFormatter: sentimentindicator1 //backgroundColor 
      valueColorFormatter: sentimentindicator1text //textColors
      fontSize: medium
    }

    view metric #colorcoding_5pt {
      backgroundColorFormatter: sentimentindicator_bg_5pt //backgroundColor 
      valueColorFormatter: sentimentindicator_text_5pt //textColors
      fontSize: medium
    }

    view metric #viewnpssegment {
      backgroundColorFormatter: sentimentindicator2a //backgroundColor 
      valueColorFormatter: sentimentindicator2text //textColors
      fontSize: medium
    }

    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext2
      backgroundColorFormatter: sentimentindicator2
      fontSize: medium
    }

    group question {
      label: "All Comments"
      comment: textAnalyticsDataset_Dining.overallScore:text
      filter expression #excludeBlankResponses {
        value: textAnalyticsDataset_Dining.overallScore:text != ""
      }
    }
    column response #comments {
      header: "Location: " + surveyDataset_TA:LocationName
      footer: @reportConfig.intvdate_ta
      view: viewComments
      enableColumnFilter: true
    }
    column value #valueColumn_OpenEnds {
      label: "Comment Field"
      value: textAnalyticsDataset_Dining.overallScore:variable
      enableColumnFilter: true
      width: 125px
    }

    column value #LocationName {
      label: "Location"
      value: surveyDataset_TA:LocationName
      enableColumnFilter: true
      //value: surveyDataset:SitesHierarchy
      width: 125px
    }

    column value #StoreName {
      label: "Store / Restaurant"
      value: surveyDataset_TA:STORE_INFO
      enableColumnFilter: true
      //value: surveyDataset_TA:SitesHierarchy
      width: 125px
    }

    column metric #metricColumn_overall_sentiment {
      label: "Overall Sentiment"
      value: score(textAnalyticsDataset_Dining:PosNegNeutralGroupsOverallSentiment)
      //value: textAnalyticsDataset_Dining:overallAverageTASet1()
      view: sentimentperformance
      format: sentimentindicatortextValue2
      enableColumnFilter: true
      width: 150px
    }


    column metric #metricColumn_NPSSegment {
      label: "NPS® Segment"
      value: score(surveyDataset_TA:NPSVal)
      format: npssegmentindicatortextValue2
      target: 3
      view: viewnpssegment
      width: 120px
      align: center
      enableColumnFilter: true

    }

    // column metric #metricColumn_NPS {
    //   label: "NPS"
    //   value: score(@reportConfig.nps_qid_ta)
    //   enableColumnFilter: true
    //   //filterable: true
    //   width: 125px
    //   align: center
    //   view: colorcoding


    // }

    // column metric #metricColumn_OSAT {
    //   label: "SAT"
    //   value: score(@reportConfig.osat_qid_ta)
    //   enableColumnFilter: true
    //   width: 125px
    //   align: center
    //   view: colorcoding_5pt
    // }

    // column metric #metricColumn_Value {
    //   label: "Value"
    //   value: score(@reportConfig.value_qid_ta)
    //   enableColumnFilter: true
    //   width: 125px
    //   align: center
    //   view: colorcoding_5pt
    // }

    view comment #viewComments {
      lines: 10
    }

  } // end widget
} // end page