//https://pr.staging.firmglobal.net/apps/editor/191375/page_133
title "MEMBER JOURNEY DEMO"

config editor {
  trace: true
}

config hub {
  hub: 579




  dataset survey #surveyDataset_Combo {
    publicName: p291026315346
    variable singleChoice #OA2__NPS {
      table: surveyDataset_Combo:
      value: recode(surveyDataset_Combo:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_Combo:
      value: recode(surveyDataset_Combo:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_Combo {
      table: surveyDataset_Combo:
      value: iif(selected(surveyDataset_Combo:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_Combo:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_Combo:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }

  dataset survey #surveyDataset_NP {
    publicName: p931921245712
    variable singleChoice #NP_ACR1 {
      label: "Availability of primary care doctors in network"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_AC1
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_ACR2 {
      label: "Availability of specialist doctors in network"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_AC2
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_ACR3 {
      label: "Availability of labs/testing sites in network"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_AC3
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_ACR4 {
      label: "Availability of pharmacies that accept your plan"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_AC4
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_BCR1 {
      label: "Coverage of doctor visits"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_BC1
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_BCR2 {
      label: "Coverage of labs/tests"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_BC2
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_BCR3 {
      label: "Value of benefits"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_BC3
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_PXR1 {
      label: "Ease of obtaining prescriptions"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_PX1
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_PXR2 {
      label: "Cost of prescriptions"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_PX2
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_PXR3 {
      label: "Coverage of prescribed medications"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_PX3
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_UPR1 {
      label: "Ease of getting benefits information"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_UP1
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_UPR2 {
      label: "Ease of getting provider information"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_UP2
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_UPR3 {
      label: "Wellness plan"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_UP3
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_UPR4 {
      label: "Plan rep's response to questions"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_UP4
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_UPR5 {
      label: "Ease of submitting claim"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_UP5
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_UPR6 {
      label: "Timeliness of claim reimbursement"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_UP6
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_YHR1 {
      label: "Understand your responsibilites in care"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_YH1
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_YHR2 {
      label: "Know what you can do to affect health"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_YH2
      option code {
        code: "1"
        score: 0
        label: "Very Poor"
      }
      option code {
        code: "2"
        score: 25
        label: "Poor"
      }
      option code {
        code: "3"
        score: 50
        label: "Fair"
      }
      option code {
        code: "4"
        score: 75
        label: "Good"
      }
      option code {
        code: "5"
        score: 100
        label: "Very Good"
      }
    }
    variable singleChoice #NP_BIR1 {
      label: "Health plan is a market leader"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_BI1
      option code {
        code: "1"
        score: 0
        label: "Completely disagree"
      }
      option code {
        code: "2"
        score: 25
        label: "Somewhat disagree"
      }
      option code {
        code: "3"
        score: 50
        label: "Neither agree nor disagree"
      }
      option code {
        code: "4"
        score: 75
        label: "Somewhat agree"
      }
      option code {
        code: "5"
        score: 100
        label: "Completely agree"
      }
    }
    variable singleChoice #NP_BIR2 {
      label: "Health plan is trustworthy"
      table: surveyDataset_NP:
      value: surveyDataset_NP:NP_BI2
      option code {
        code: "1"
        score: 0
        label: "Completely disagree"
      }
      option code {
        code: "2"
        score: 25
        label: "Somewhat disagree"
      }
      option code {
        code: "3"
        score: 50
        label: "Neither agree nor disagree"
      }
      option code {
        code: "4"
        score: 75
        label: "Somewhat agree"
      }
      option code {
        code: "5"
        score: 100
        label: "Completely agree"
      }
    }
    variable grid #AccessToCareGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_ACR1, surveyDataset_NP:NP_ACR2, surveyDataset_NP:NP_ACR3, surveyDataset_NP:NP_ACR4)
    }
    variable grid #BenefitsCoverageGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_BCR1, surveyDataset_NP:NP_BCR2, surveyDataset_NP:NP_BCR3)
    }
    variable grid #PrescriptionsGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_PXR1, surveyDataset_NP:NP_PXR2, surveyDataset_NP:NP_PXR3)
    }
    variable grid #UsingHPGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_UPR1, surveyDataset_NP:NP_UPR2, surveyDataset_NP:NP_UPR3, surveyDataset_NP:NP_UPR4, surveyDataset_NP:NP_UPR5, surveyDataset_NP:NP_UPR6)
    }
    variable grid #YourHealthGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_YHR1, surveyDataset_NP:NP_YHR2)
    }
    variable grid #BrandImageGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_BIR1, surveyDataset_NP:NP_BIR2)
    }
    variable grid #DoctorsGrid {
      table: surveyDataset_NP:
      value: vlist(surveyDataset_NP:NP_DR2, surveyDataset_NP:NP_DR4)
    }
    variable singleChoice #OA2__NPS {
      table: surveyDataset_NP:
      value: recode(surveyDataset_NP:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_NP:
      value: recode(surveyDataset_NP:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_NP {
      table: surveyDataset_NP:
      value: iif(selected(surveyDataset_NP:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_NP:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_NP:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  vtable split #AccessToCare {
    source: surveyDataset_NP:AccessToCareGrid
  }
  vtable split #BenefitsCoverage {
    source: surveyDataset_NP:BenefitsCoverageGrid
  }
  vtable split #Prescriptions {
    source: surveyDataset_NP:PrescriptionsGrid
  }
  vtable split #UsingHP {
    source: surveyDataset_NP:UsingHPGrid
  }
  vtable split #YourHealth {
    source: surveyDataset_NP:YourHealthGrid
  }
  vtable split #BrandImage {
    source: surveyDataset_NP:BrandImageGrid
  }
  vtable split #Doctors {
    source: surveyDataset_NP:DoctorsGrid
  }
  variable auto #Dial__gridTile_1__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_AC1, surveyDataset_NP:NP_AC2, surveyDataset_NP:NP_AC3, surveyDataset_NP:NP_AC4)
  }
  variable auto #Dial__gridTile_2__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_BC1, surveyDataset_NP:NP_BC2, surveyDataset_NP:NP_BC3)
  }
  variable auto #Dial__gridTile_3__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_PX1, surveyDataset_NP:NP_PX2, surveyDataset_NP:NP_PX3)
  }
  variable auto #Dial__gridTile_4__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_UP1, surveyDataset_NP:NP_UP2, surveyDataset_NP:NP_UP3, surveyDataset_NP:NP_UP4, surveyDataset_NP:NP_UP5, surveyDataset_NP:NP_UP6)
  }
  variable auto #Dial__gridTile_5__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_YH1, surveyDataset_NP:NP_YH2)
  }
  variable auto #Dial__gridTile_6__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_BI1, surveyDataset_NP:NP_BI2)
  }
  variable auto #Dial__gridTile_7__variable {
    table: surveyDataset_NP:
    value: VList(surveyDataset_NP:NP_DR2, surveyDataset_NP:NP_DR4)
  }

  dataset survey #surveyDataset_SA {
    publicName: p328843140028
    variable grid #ProviderAvailabilityGrid {
      table: surveyDataset_SA:
      value: vlist(surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8)
    }
    variable grid #RxAvailabilityGrid {
      table: surveyDataset_SA:
      value: vlist(surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4, surveyDataset_SA:SA_RX5)
    }
    variable grid #PremiumCoveragesGrid {
      table: surveyDataset_SA:
      value: vlist(surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3)
    }
    variable singleChoice #OA2__NPS {
      table: surveyDataset_SA:
      value: recode(surveyDataset_SA:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_SA:
      value: recode(surveyDataset_SA:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_SA {
      table: surveyDataset_SA:
      value: iif(selected(surveyDataset_SA:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_SA:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_SA:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  vtable split #ProviderAvailability {
    source: surveyDataset_SA:ProviderAvailabilityGrid
  }
  vtable split #RxAvailability {
    source: surveyDataset_SA:RxAvailabilityGrid
  }
  vtable split #PremiumCoverages {
    source: surveyDataset_SA:PremiumCoveragesGrid
  }
  variable auto #Dial__gridTile_8__variable {
    table: surveyDataset_SA:
    value: VList(surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8)
  }
  variable auto #Dial__gridTile_9__variable {
    table: surveyDataset_SA:
    value: VList(surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4, surveyDataset_SA:SA_RX5)
  }
  variable auto #Dial__gridTile_10__variable {
    table: surveyDataset_SA:
    value: VList(surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3)
  }
  variable auto #Dial__gridTile_11__variable {
    table: surveyDataset_SA:
    value: VList(surveyDataset_SA:SA_SB1)
  }

  dataset survey #surveyDataset_EN {
    publicName: p132177326256
  }

  dataset survey #surveyDataset_SO {
    publicName: p700259985250
  }

  dataset survey #surveyDataset_PT {
    publicName: p951947950682
  }

  dataset survey #surveyDataset_CO {
    publicName: p393201032957
  }

  dataset survey #surveyDataset_FC {
    publicName: p588253035121
  }

  dataset survey #surveyDataset_AC {
    publicName: p417223780420
    variable grid #MakingApptsGrid {
      table: surveyDataset_AC:
      value: vlist(surveyDataset_AC:AC_MA2, surveyDataset_AC:AC_MA3, surveyDataset_AC:AC_MA4)
    }
    variable singleChoice #OA2__NPS {
      table: surveyDataset_AC:
      value: recode(surveyDataset_AC:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_AC:
      value: recode(surveyDataset_AC:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_AC {
      table: surveyDataset_AC:
      value: iif(selected(surveyDataset_AC:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_AC:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_AC:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  vtable split #MakingAppts {
    source: surveyDataset_AC:MakingApptsGrid
  }
  variable auto #Dial__gridTile_22__variable {
    table: surveyDataset_AC:
    value: VList(surveyDataset_AC:AC_MA2, surveyDataset_AC:AC_MA3, surveyDataset_AC:AC_MA4)
  }

  dataset survey #surveyDataset_MP {
    publicName: p364207198558
  }

  dataset survey #surveyDataset_CR {
    publicName: p193236180368
  }

  dataset survey #surveyDataset_CM {
    publicName: p887894748791
  }

  dataset survey #surveyDataset_SB {
    publicName: p110556283834
  }

  dataset survey #surveyDataset_RXCombo {
    publicName: p779568282910
    variable singleChoice #OA2__NPS {
      table: surveyDataset_Combo:
      value: recode(surveyDataset_RXCombo:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_RXCombo:
      value: recode(surveyDataset_RXCombo:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_RXCombo {
      table: surveyDataset_Combo:
      value: iif(selected(surveyDataset_RXCombo:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_RXCombo:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_RXCombo:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  dataset survey #surveyDataset_RP {
    publicName: p333859452405
    variable grid #RXPreAuthGrid {
      table: surveyDataset_RP:
      value: vlist(surveyDataset_RP:RP_PA3, surveyDataset_RP:RP_PA6)
    }
    variable singleChoice #OA2__NPS {
      table: surveyDataset_RP:
      value: recode(surveyDataset_RP:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_RP:
      value: recode(surveyDataset_RP:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_RP {
      table: surveyDataset_RP:
      value: iif(selected(surveyDataset_RP:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_RP:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_RP:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  vtable split #RXPreAuth {
    source: surveyDataset_RP:RXPreAuthGrid
  }
  variable auto #Dial__gridTile_32__variable {
    table: surveyDataset_RP:
    value: VList(surveyDataset_RP:RP_PA3, surveyDataset_RP:RP_PA6)
  }

  dataset survey #surveyDataset_GP {
    publicName: p538182290991
    variable grid #RetailRXGrid {
      table: surveyDataset_GP:
      value: vlist(surveyDataset_GP:GP_RX2, surveyDataset_GP:GP_RX3, surveyDataset_GP:GP_RX4, surveyDataset_GP:GP_RX5, surveyDataset_GP:GP_RX6)
    }
    variable grid #MailRXGrid {
      table: surveyDataset_GP:
      value: vlist(surveyDataset_GP:GP_MX2, surveyDataset_GP:GP_MX3, surveyDataset_GP:GP_MX4, surveyDataset_GP:GP_MX5, surveyDataset_GP:GP_MX6)
    }
    variable singleChoice #OA2__NPS {
      table: surveyDataset_GP:
      value: recode(surveyDataset_GP:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_GP:
      value: recode(surveyDataset_GP:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_GP {
      table: surveyDataset_GP:
      value: iif(selected(surveyDataset_GP:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_GP:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_GP:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  vtable split #RetailRX {
    source: surveyDataset_GP:RetailRXGrid
  }
  vtable split #MailRX {
    source: surveyDataset_GP:MailRXGrid
  }
  variable auto #Dial__gridTile_33__variable {
    table: surveyDataset_GP:
    value: VList(surveyDataset_GP:GP_RX2, surveyDataset_GP:GP_RX3, surveyDataset_GP:GP_RX4, surveyDataset_GP:GP_RX5, surveyDataset_GP:GP_RX6)
  }
  variable auto #Dial__gridTile_34__variable {
    table: surveyDataset_GP:
    value: VList(surveyDataset_GP:GP_MX2, surveyDataset_GP:GP_MX3, surveyDataset_GP:GP_MX4, surveyDataset_GP:GP_MX5, surveyDataset_GP:GP_MX6)
  }

  dataset survey #surveyDataset_CX {
    publicName: p543363096658
    variable grid #ConRXGrid {
      table: surveyDataset_CX:
      value: vlist(surveyDataset_CX:CX_CS2, surveyDataset_CX:CX_CS3, surveyDataset_CX:CX_CS4)
    }
    variable singleChoice #OA2__NPS {
      table: surveyDataset_CX:
      value: recode(surveyDataset_CX:OA2, @_NPS)
      label: "NPS"
    }
    variable singleChoice #OA2__scale10To3 {
      table: surveyDataset_CX:
      value: recode(surveyDataset_CX:OA2, @_scale10To3)
      label: "NPS"
    }
    variable singleChoice #NPSRecode_CX {
      table: surveyDataset_CX:
      value: iif(selected(surveyDataset_CX:OA2, "0", "1", "2", "3", "4", "5", "6"), "Detractor", iif(selected(surveyDataset_CX:OA2, "7", "8"), "Passive", iif(selected(surveyDataset_CX:OA2, "9", "10"), "Promoter")))
      option code {
        code: "Promoter"
        label: "Promoter"
      }
      option code {
        code: "Passive"
        label: "Passive"
      }
      option code {
        code: "Detractor"
        label: "Detractor"
      }
    }
  }
  vtable split #ConRX {
    source: surveyDataset_CX:ConRXGrid
  }
  variable auto #Dial__gridTile_35__variable {
    table: surveyDataset_CX:
    value: VList(surveyDataset_CX:CX_CS2, surveyDataset_CX:CX_CS3, surveyDataset_CX:CX_CS4)
  }

  dataset survey #surveyDataset_CS {
    publicName: p394814974667
  }

  dataset survey #surveyDataset_MC {
    publicName: p107001804067
  }

  dataset survey #surveyDataset_XC {
    publicName: p929431604982
  }

  dataset survey #surveyDataset_SC {
    publicName: p559326564531
  }

  dataset survey #surveyDataset_RC {
    publicName: p102973223258
  }

  dataset survey #surveyDataset_DI {
    publicName: p857124398263
  }

  dataset cases #cases {
    publicName: am
  }



  variableSet #variableSet_NP {
    label: "Selector"
    table: surveyDataset_NP:
    variables: surveyDataset_NP:ITLOB, surveyDataset_NP:ITGENDER, surveyDataset_NP:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_NP:ITLOB
    }
  }
  variableSet #variableSet_SA {
    label: "Selector"
    table: surveyDataset_SA:
    variables: surveyDataset_SA:ITLOB, surveyDataset_SA:ITGENDER, surveyDataset_SA:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_SA:ITLOB
    }
  }
  variableSet #variableSet_AC {
    label: "Selector"
    table: surveyDataset_AC:
    variables: surveyDataset_AC:ITLOB, surveyDataset_AC:ITGENDER, surveyDataset_AC:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_AC:ITLOB
    }
  }
  variableSet #variableSet_RXCombo {
    label: "Selector"
    table: surveyDataset_RXCombo:
    variables: surveyDataset_RXCombo:ITLOB, surveyDataset_RXCombo:ITGENDER, surveyDataset_RXCombo:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_RXCombo:ITLOB
    }
  }
  variableSet #variableSet_RP {
    label: "Selector"
    table: surveyDataset_RP:
    variables: surveyDataset_RP:ITLOB, surveyDataset_RP:ITGENDER, surveyDataset_RP:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_RP:ITLOB
    }
  }
  variableSet #variableSet_GP {
    label: "Selector"
    table: surveyDataset_GP:
    variables: surveyDataset_GP:ITLOB, surveyDataset_GP:ITGENDER, surveyDataset_GP:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_GP:ITLOB
    }
  }
  variableSet #variableSet_CX {
    label: "Selector"
    table: surveyDataset_CX:
    variables: surveyDataset_CX:ITLOB, surveyDataset_CX:ITGENDER, surveyDataset_CX:ITMEMST
    hint visualDesigner #selectHint {
      defaultOption: surveyDataset_CX:ITLOB
    }
  }
}
custom properties #operationalProperties {
  combo: surveyDataset_Combo:combined_sourceid = "p291026315346"
  foundations: surveyDataset_Combo:combined_sourceid = "p931921245712"
  sales: surveyDataset_Combo:combined_sourceid = "p328843140028"
  accesstocare: surveyDataset_Combo:combined_sourceid = "p417223780420"
  rxmgmt: surveyDataset_Combo:combined_sourceid = "p779568282910"
  rxpreauth: surveyDataset_Combo:combined_sourceid = "p333859452405"
  gettingrx: surveyDataset_Combo:combined_sourceid = "p538182290991"
  conrx: surveyDataset_Combo:combined_sourceid = "p543363096658"
}
config queryOptions {
  // added automatically during report creation
  boolNullsAsFalse: false
  explicitLevelAggregation: true
}

layoutArea toolbar {
  useDynamicFilters: true
  filter reportingPeriod #reportingPeriodFilter {
    label: "Time Period"
  }
  filter multiselect #fromQuestionFilter_Combo_LOB {
    optionsFrom: surveyDataset_Combo:ITLOB
    label: "Line of Business"
  }
  filter multiselect #fromQuestionFilter_Combo_PLAN {
    optionsFrom: surveyDataset_Combo:ITPLAN_TY
    label: "Plan Type"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_Combo_CONTRACT {
    optionsFrom: surveyDataset_Combo:ITH_CONTRACT
    label: "Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_Combo_GENDER {
    optionsFrom: surveyDataset_Combo:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "Gender"
  }
  filter multiselect #fromQuestionFilter_Combo_RACE {
    optionsFrom: surveyDataset_Combo:ITRACE
    label: "Race"
  }
  filter multiselect #fromQuestionFilter_Combo_MEMST {
    optionsFrom: surveyDataset_Combo:ITMEMST
    label: "Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_Combo_OA1 {
    optionsFrom: surveyDataset_Combo:OA1
  }
  filter multiselect #fromQuestionFilter_NP_LOB {
    optionsFrom: surveyDataset_NP:ITLOB
    label: "(FOUNDATIONS) Line of Business"
  }
  filter multiselect #fromQuestionFilter_NP_PLAN {
    optionsFrom: surveyDataset_NP:ITPLAN_TY
    label: "(FOUNDATIONS) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_NP_CONTRACT {
    optionsFrom: surveyDataset_NP:ITH_CONTRACT
    label: "(FOUNDATIONS) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_NP_GENDER {
    optionsFrom: surveyDataset_NP:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(FOUNDATIONS) Gender"
  }
  filter multiselect #fromQuestionFilter_NP_RACE {
    optionsFrom: surveyDataset_NP:ITRACE
    label: "(FOUNDATIONS) Race"
  }
  filter multiselect #fromQuestionFilter_NP_MEMST {
    optionsFrom: surveyDataset_NP:ITMEMST
    label: "(FOUNDATIONS) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_SA_LOB {
    optionsFrom: surveyDataset_SA:ITLOB
    label: "(SALES) Line of Business"
  }
  filter multiselect #fromQuestionFilter_SA_PLAN {
    optionsFrom: surveyDataset_SA:ITPLAN_TY
    label: "(SALES) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_SA_CONTRACT {
    optionsFrom: surveyDataset_SA:ITH_CONTRACT
    label: "(SALES) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_SA_GENDER {
    optionsFrom: surveyDataset_SA:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(SALES) Gender"
  }
  filter multiselect #fromQuestionFilter_SA_RACE {
    optionsFrom: surveyDataset_SA:ITRACE
    label: "(SALES) Race"
  }
  filter multiselect #fromQuestionFilter_SA_MEMST {
    optionsFrom: surveyDataset_SA:ITMEMST
    label: "(SALES) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_SA_OA1 {
    optionsFrom: surveyDataset_SA:OA1
    label: "(SALES) Overall Experience"
  }
  filter multiselect #fromQuestionFilter_AC_LOB {
    optionsFrom: surveyDataset_AC:ITLOB
    label: "(ACCESS TO CARE) Line of Business"
  }
  filter multiselect #fromQuestionFilter_AC_PLAN {
    optionsFrom: surveyDataset_AC:ITPLAN_TY
    label: "(ACCESS TO CARE) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_AC_CONTRACT {
    optionsFrom: surveyDataset_AC:ITH_CONTRACT
    label: "(ACCESS TO CARE) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_AC_GENDER {
    optionsFrom: surveyDataset_AC:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(ACCESS TO CARE) Gender"
  }
  filter multiselect #fromQuestionFilter_AC_RACE {
    optionsFrom: surveyDataset_AC:ITRACE
    label: "(ACCESS TO CARE) Race"
  }
  filter multiselect #fromQuestionFilter_AC_MEMST {
    optionsFrom: surveyDataset_AC:ITMEMST
    label: "(ACCESS TO CARE) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_AC_OA1 {
    optionsFrom: surveyDataset_AC:OA1
    label: "(ACCESS TO CARE) Overall Experience"
  }
  filter singleselect #fromQuestionFilter_AC_MA1 {
    optionsFrom: surveyDataset_AC:AC_MA1
    label: "(ACCESS TO CARE) Type of care needed"
  }
  filter multiselect #fromQuestionFilter_RXCombo_LOB {
    optionsFrom: surveyDataset_RXCombo:ITLOB
    label: "(RX MGMT) Line of Business"
  }
  filter multiselect #fromQuestionFilter_RXCombo_PLAN {
    optionsFrom: surveyDataset_RXCombo:ITPLAN_TY
    label: "(RX MGMT) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_RXCombo_CONTRACT {
    optionsFrom: surveyDataset_RXCombo:ITH_CONTRACT
    label: "(RX MGMT) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_RXCombo_GENDER {
    optionsFrom: surveyDataset_RXCombo:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(RX MGMT) Gender"
  }
  filter multiselect #fromQuestionFilter_RXCombo_RACE {
    optionsFrom: surveyDataset_RXCombo:ITRACE
    label: "(RX MGMT) Race"
  }
  filter multiselect #fromQuestionFilter_RXCombo_MEMST {
    optionsFrom: surveyDataset_RXCombo:ITMEMST
    label: "(RX MGMT) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_RXCombo_OA1 {
    optionsFrom: surveyDataset_RXCombo:OA1
    label: "(RX MGMT) Overall Experience"
  }
  filter multiselect #fromQuestionFilter_RP_LOB {
    optionsFrom: surveyDataset_RP:ITLOB
    label: "(RX PREAUTH) Line of Business"
  }
  filter multiselect #fromQuestionFilter_RP_PLAN {
    optionsFrom: surveyDataset_RP:ITPLAN_TY
    label: "(RX PREAUTH) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_RP_CONTRACT {
    optionsFrom: surveyDataset_RP:ITH_CONTRACT
    label: "(RX PREAUTH) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_RP_GENDER {
    optionsFrom: surveyDataset_RP:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(RX PREAUTH) Gender"
  }
  filter multiselect #fromQuestionFilter_RP_RACE {
    optionsFrom: surveyDataset_RP:ITRACE
    label: "(RX PREAUTH) Race"
  }
  filter multiselect #fromQuestionFilter_RP_MEMST {
    optionsFrom: surveyDataset_RP:ITMEMST
    label: "(RX PREAUTH) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_RP_OA1 {
    optionsFrom: surveyDataset_RP:OA1
    label: "(RX PREAUTH) Overall Experience"
  }
  filter singleselect #fromQuestionFilter_RP_PA4 {
    optionsFrom: surveyDataset_RP:RP_PA4
    label: "(RX PREAUTH) Preauthorization was denied"
  }
  filter multiselect #fromQuestionFilter_GP_LOB {
    optionsFrom: surveyDataset_GP:ITLOB
    label: "(GETTING RX) Line of Business"
  }
  filter multiselect #fromQuestionFilter_GP_PLAN {
    optionsFrom: surveyDataset_GP:ITPLAN_TY
    label: "(GETTING RX) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_GP_CONTRACT {
    optionsFrom: surveyDataset_GP:ITH_CONTRACT
    label: "(GETTING RX) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_GP_GENDER {
    optionsFrom: surveyDataset_GP:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(GETTING RX) Gender"
  }
  filter multiselect #fromQuestionFilter_GP_RACE {
    optionsFrom: surveyDataset_GP:ITRACE
    label: "(GETTING RX) Race"
  }
  filter multiselect #fromQuestionFilter_GP_MEMST {
    optionsFrom: surveyDataset_GP:ITMEMST
    label: "(GETTING RX) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_GP_OA1 {
    optionsFrom: surveyDataset_GP:OA1
    label: "(GETTING RX) Overall Experience"
  }
  filter multiselect #fromQuestionFilter_CX_LOB {
    optionsFrom: surveyDataset_CX:ITLOB
    label: "(CON RX) Line of Business"
  }
  filter multiselect #fromQuestionFilter_CX_PLAN {
    optionsFrom: surveyDataset_CX:ITPLAN_TY
    label: "(CON RX) Plan Type "
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_CX_CONTRACT {
    optionsFrom: surveyDataset_CX:ITH_CONTRACT
    label: "(CON RX) Contract"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_CX_GENDER {
    optionsFrom: surveyDataset_CX:ITGENDER
    sortOrder: "ascending"
    hide: false
    label: "(CON RX) Gender"
  }
  filter multiselect #fromQuestionFilter_CX_RACE {
    optionsFrom: surveyDataset_GP:ITRACE
    label: "(CON RX) Race"
  }
  filter multiselect #fromQuestionFilter_CX_MEMST {
    optionsFrom: surveyDataset_CX:ITMEMST
    label: "(CON RX) Member State"
    sortOrder: "ascending"
  }
  filter multiselect #fromQuestionFilter_CX_OA1 {
    optionsFrom: surveyDataset_CX:OA1
    label: "(CON RX) Overall Experience"
  }
}

config style #styleConfig {
  theme: "modern"
}

config pdfExport {
  pageSize: "Letter"
  pageOrientation: "landscape", "portrait"
  pageScaling: fitToWidth
  exportMode: htmlToPdf
  version: 2
  allowFileNaming: true
  pageMargins: 0.4
}

config headerBarTheme {
  headerBackgroundColor: ""
  headerBottomLineColor: ""
  tabsBackgroundColor: ""
  tabsTextColor: ""
  activeTabColor: #2b3584
}

config calendarOptions #calendarOptionsConfig {
  weekRule: "firstDay"
}

config mobile {
  showShareButton: true
}

config report #reportConfig {
  logo: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Logos/PG_Logo_RGB_Navy.png"
  formatter number #n_EqualsWithComma_baseFormatter {
    label: "base, formatter"
    prefix: "(n="
    numberDecimals: 0
    postfix: ")"
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
  }

  formatter number #N_Equals_baseFormatter {
    label: "Base formatter"
    prefix: "(N="
    numberDecimals: 0
    postfix: ")"
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
  }

  formatter date #dateDefaultFormat {
    formatString: "MMM DD YYYY"
    emptyValue: " "
  }

  formatter period #weekFormat {
    inputFormat: "YYYYWW"
    formatString: "{start:MMM DD YYYY}"
    datePart: calendarWeek
  }

  formatter color #kpiColorDefaultFormatter {
    label: "Red Amber Green Percent (KPI)-2"
    thresholds: #12A1A1 > 75, #4B82F0 > 50, #E27508 > 25, #D02541 <= 25
    defaultValue: #ffffff = 0
  }
  formatter color #SurveyResponseColorScaledMeanScoreFormatter {
    label: "Red Amber Green Scaled Mean"
    thresholds: #12A1A1 > 75, #4B82F0 > 50, #E27508 > 25, #D02541 <= 25
  }
  formatter color #SurveyResponseColorPastelBackgroundFormatter {
    label: "Red Amber Green Scaled Mean Background"
    thresholds: #DBFBFB > 75, #DFE9FD > 50, #FDE7D0 > 25, #F9DBE0 <= 25
  }
  formatter color #gridDefaultBackgroundColorFormatter {
    label: "Red Amber Green Background"
    thresholds: #D3EFDA >= 95%, #FFFFE0 >= 90%, #F7D4D4 < 90%
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter color #DifferenceBlackRedFormatter {
    label: "Black Red Numeric base"
    thresholds: #000000 >= 30, #D02525 < 30
  }
  formatter color #colorFormatter_Promoters {
    thresholds: #519B14 >= 0, #519B14 < 100%
    label: "Promoters Color"
  }
  formatter color #colorFormatter_Passives {
    thresholds: #FF6D00 >= 0, #FF6D00 < 100%
    label: "Passives Color"
  }
  formatter color #colorFormatter_Detractors {
    thresholds: #FA5263 >= 0, #FA5263 < 100%
    label: "Detractors Color"
  }
  palette #NPSColorPalette {
    label: "NPS Color Palette"
    colors: "#FA5263", "#FF6D00", "#519B14"
  }
  palette #Single_Red_Color_Bar {
    label: "Single Red Color Bar"
    colors: "#D02541"
  }

  formatter number #NoDecimalsNumberFormatter {
    label: "No Decimals"
    numberDecimals: 0
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
    emptyValue: "-"
  }
  formatter number #OneDecimalNumberFormatter {
    label: "One Decimal"
    numberDecimals: 1
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: true
    ordinal: false
    emptyValue: "-"
  }
  formatter number #percentNoDecimalDefaultFormatter {
    label: "Percent No Decimal"
    numberDecimals: 0
    postfix: "%"
    emptyValue: "-"
    prefix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
  }
  formatter number #percentScaleNoDecimalDefaultFormatter {
    label: "Percent No Decimal Scale"
    numberDecimals: 0
    postfix: "%"
    emptyValue: "-"
    prefix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
  }
  formatter number #PercentOneDecimalFormatter {
    label: "Percent One Decimal"
    postfix: "%"
    emptyValue: "-"
    prefix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: true
    ordinal: false
    numberDecimals: 1
  }
  formatter number #numberFormatter {
    decimalSeparator: "."
    integerSeparator: ","
  }
  formatter number #bigNumberFormatter {
    label: "No Decimals"
    numberDecimals: 0
    prefix: ""
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter number #bigNumberScaleFormatter {
    label: "No Decimals Scale"
    numberDecimals: 0
    prefix: ""
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter number #floatDefaultFormatter {
    label: "Two Decimals with No Empty Value"
    numberDecimals: 2
    prefix: ""
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter number #percentNoDecimal {
    label: "Percent No Decimal"
    numberDecimals: 0
    postfix: "%"
    emptyValue: "-"
    prefix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
// This default formatter was added to CDL when it was overridden in the widget library
  }
  formatter number #baseDefaultFormatter {
    label: "Base formatter"
    prefix: "(N="
    numberDecimals: 0
    postfix: ")"
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
// This default formatter was added to CDL when it was overridden in the widget library
  }
}





page #page_133 {
  label: "MEMBER JOURNEY"
  widget canvas #canvasWidget {
    label: "Canvas"
    container: container position {
      width: 1368px
      height: 800px
      background: "url('/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Moments%20that%20matter%20Dashboard_Fan.png') 0% 0% / cover no-repeat"
      area #area {
        position: "absolute"
        top: "444px"
        left: "467px"
      }
      area #area_2 {
        position: "absolute"
        top: "454px"
        left: "771px"
      }
      area #area_3 {
        position: "absolute"
        top: "352px"
        left: "1105px"
      }
      area #area_4 {
        position: "absolute"
        top: "508px"
        left: "27px"
      }
      area #area_5 {
        position: "absolute"
        top: "215px"
        left: "1019px"
      }
      area #area_6 {
        position: "absolute"
        top: "81px"
        left: "869px"
      }
      area #area_7 {
        position: "absolute"
        top: "520px"
        left: "1120px"
      }
      area #area_8 {
        position: "absolute"
        top: "17px"
        left: "686px"
      }
      area #area_9 {
        position: "absolute"
        top: "349px"
        left: "82px"
      }
      area #area_10 {
        position: "absolute"
        top: "192px"
        left: "164px"
      }
      area #area_11 {
        position: "absolute"
        top: "78px"
        left: "295px"
      }
      area #area_12 {
        position: "absolute"
        top: "20px"
        left: "486px"
      }
      area #area_14 {
        position: "absolute"
        top: "486px"
        left: "215px"
      }
      area #area_15 {
        position: "absolute"
        top: "353px"
        left: "264px"
      }
      area #area_16 {
        position: "absolute"
        top: "259px"
        left: "381px"
      }
      area #area_17 {
        position: "absolute"
        top: "176px"
        left: "530px"
      }
      area #area_18 {
        position: "absolute"
        top: "611px"
        left: "1042px"
      }
      area #area_19 {
        position: "absolute"
        top: "473px"
        left: "1008px"
      }
      area #area_22 {
        position: "absolute"
        top: "178px"
        left: "703px"
      }
      area #area_20 {
        position: "absolute"
        top: "497px"
        left: "1041px"
      }
      area #area_21 {
        position: "absolute"
        top: "599px"
        left: "210px"
      }
      area #area_23 {
        position: "absolute"
        top: "175px"
        left: "703px"
      }
      area #area_24 {
        position: "absolute"
        top: "241px"
        left: "838px"
      }
      area #area_25 {
        position: "absolute"
        top: "338px"
        left: "996px"
      }
      area #area_26 {
        top: "599px"
        left: "335px"
        position: "absolute"
      }
      area #area_27 {
        position: "absolute"
        top: "508px"
        left: "364px"
      }
      area #area_28 {
        position: "absolute"
        top: "425px"
        left: "403px"
      }
      area #area_29 {
        position: "absolute"
        top: "352px"
        left: "495px"
      }
      area #area_30 {
        position: "absolute"
        top: "334px"
        left: "586px"
      }
      area #area_31 {
        position: "absolute"
        top: "355px"
        left: "713px"
      }
    }
    cardTransparent: true
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/people_business_consumer-15.png"
      areaId: "area"
      style #style {
        width: "159px"
      }
    }
    tile image #imageTile_2 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/people_business_consumer-16.png"
      areaId: "area_2"
      style #style {
        width: "152px"
      }
    }
    tile image #imageTile_3 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-13.png"
      areaId: "area_3"
      style #style {
        width: 200px
      }
      label: "Recommend_Care"
    }
    tile image #imageTile_4 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-04.png"
      areaId: "area_4"
      style #style {
        width: "200px"
      }
      label: "Sales"
    }
    tile image #imageTile_5 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-12.png"
      areaId: "area_5"
      style #style {
        width: 200px
      }
      label: "Costs"
    }
    tile image #imageTile_6 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-10.png"
      areaId: "area_6"
      style #style {
        width: 200px
      }
      label: "Customer_Service"
    }
    tile image #imageTile_7 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-11.png"
      areaId: "area_7"
      style #style {
        width: 200px
      }
      label: "Disenrollement"
    }
    tile image #imageTile_8 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-09.png"
      areaId: "area_8"
      style #style {
        width: 200px
      }
      label: "Rx_Management"
    }
    tile image #imageTile_9 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-05.png"
      areaId: "area_9"
      style #style {
        width: 200px
      }
      label: "Enrollement"
    }
    tile image #imageTile_10 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-06.png"
      areaId: "area_10"
      style #style {
        width: 200px
      }
      label: "Onboarding"
    }
    tile image #imageTile_11 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-07.png"
      areaId: "area_11"
      style #style {
        width: 200px
      }
      label: "Finding_Care"
    }
    tile image #imageTile_12 {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Demo%20File/Member%20Journey%20WIP/Moments%20that%20matter%20Dashboard_icons-08.png"
      areaId: "area_12"
      style #style {
        width: 200px
      }
      label: "Benefit_Usage"
    }
    tile text #textTile_2 {
      value: "Enrollment"
      areaId: "area_14"
      style #style {
        fontSize: 24
        color: #4b1bcd
        fontWeight: "bold"
      }
    }
    tile text #textTile_3 {
      value: "Onboarding"
      areaId: "area_15"
      style #style {
        fontSize: 24
        color: #7d5ff2
        fontWeight: "bold"
      }
    }
    tile text #textTile_4 {
      value: "Finding Care"
      areaId: "area_16"
      style #style {
        fontSize: 24
        color: #a444dd
        fontWeight: "bold"
      }
    }
    tile text #textTile_5 {
      value: "Benefit Usage"
      areaId: "area_17"
      style #style {
        fontSize: 22
        color: #ca2d76
        fontWeight: "bold"
      }
    }
    tile text #textTile_6 {
      value: "Disenrollment"
      areaId: "area_18"
      style #style {
        fontSize: 20
        color: #343e47
        fontWeight: "bold"
      }
    }
    tile text #textTile_7 {
      value: "Recommended"
      areaId: "area_19"
      style #style {
        fontSize: 24
        color: #7d868b
        fontWeight: "bold"
      }
    }
    tile text #textTile_8 {
      value: "Care"
      areaId: "area_20"
      style #style {
        fontSize: 24
        color: #7d868b
        fontWeight: "bold"
      }
    }
    tile text #textTile_9 {
      value: "Sales"
      areaId: "area_21"
      style #style {
        fontSize: 24
        color: #030862
        fontWeight: "bold"
      }
    }
    tile text #textTile_10 {
      value: "Rx Mngmnt"
      areaId: "area_23"
      style #style {
        fontSize: 24
        color: #992175
        fontWeight: "bold"
      }
    }
    tile text #textTile_11 {
      value: "Customer Service"
      areaId: "area_24"
      style #style {
        fontSize: 20
        color: #7d1773
        fontWeight: "bold"
      }
    }
    tile text #textTile_12 {
      value: "Costs"
      areaId: "area_25"
      style #style {
        fontSize: 24
        color: #540c54
        fontWeight: "bold"
      }
    }
    tile value #valueTile {
      areaId: "area_26"
      label: "NPS"
      value: 72
      style #style {
        justifyContent: "start"
        alignItems: "start"
        fontSize: 45
        color: #ffffff
        fontWeight: "bold"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_27"
      label: "NPS"
      value: 72
      style #style {
        justifyContent: "start"
        alignItems: "start"
        fontSize: 45
        color: #ffffff
        fontWeight: "bold"
      }
    }
    tile value #valueTile_3 {
      areaId: "area_28"
      label: "NPS"
      value: 72
      style #style {
        justifyContent: "start"
        alignItems: "start"
        fontSize: 45
        color: #ffffff
        fontWeight: "bold"
      }
    }
    tile value #valueTile_4 {
      areaId: "area_29"
      label: "NPS"
      value: 72
      style #style {
        justifyContent: "start"
        alignItems: "start"
        fontSize: 45
        color: #ffffff
        fontWeight: "bold"
      }
    }
    tile value #valueTile_5 {
      areaId: "area_30"
      label: "NPS"
      value: 72
      style #style {
        justifyContent: "start"
        alignItems: "start"
        fontSize: 45
        color: #ffffff
        fontWeight: "bold"
      }
    }
    tile value #valueTile_6 {
      areaId: "area_31"
      label: "NPS"
      value: 72
      style #style {
        justifyContent: "start"
        alignItems: "start"
        fontSize: 45
        color: #ffffff
        fontWeight: "bold"
      }
    }
  }
  ignoreFilters: fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1
}
page #ActionMgmt {
  label: "ACTION MANAGEMENT"
  widget caseList #caseListWidget {
    cardCorners: '20px'
    label: "Case List"
    size: "large"
    navigateTo: "ActionMgmt"
  }
  widget caseDetailsSummary #caseDetailsSummaryWidget {
    cardCorners: '20px'
    label: "Case Details Summary"
    size: "large"
    navigateTo: "ActionMgmt"
    items: "id", "name", "triggerName"
  }
  widget caseLog #caseLogWidget {
    cardCorners: '20px'
    label: "Case Log"
    size: "large"
    ignoreFiscalCalendar: true
  }
  widget caseManagement #caseManagementWidget {
    cardCorners: '20px'
    label: "Case Management"
    size: "halfwidth"
  }
  widget caseResponse #caseResponseWidget {
    cardCorners: '20px'
    label: "Case Response"
    size: "halfwidth"
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1
  config layout #layoutConfig {
    horizontalAlignmentMode: ""
  }
  hide: false
  modal: true
}











page #SA_Select_Q_by {
  label: "SA_Select_Q_by"
  widget dataGrid #dataGridWidget {
    cardCorners: '20px'
    label: "Scores by Category"
    size: medium
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_SA:ITLOB
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_SA:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_SA:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_SA:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_SA:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_SA:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_SA:OA1
          target: 77
          removeEmptyRows: true
        }
      },
      item {
        label: 'Provider Availability Composite'
        value: {
          qid: ProviderAvailability:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Existing PCP in network'
        value: {
          qid: surveyDataset_SA:SA_PA2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Existing spec in network'
        value: {
          qid: surveyDataset_SA:SA_PA4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Hospital/facility in network'
        value: {
          qid: surveyDataset_SA:SA_PA5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'PCP local'
        value: {
          qid: surveyDataset_SA:SA_PA6
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Spec local'
        value: {
          qid: surveyDataset_SA:SA_PA7
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Finding provider(s) that meet certain characteristics'
        value: {
          qid: surveyDataset_SA:SA_PA8
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Pharmacy/Rx Availability Composite'
        value: {
          qid: RxAvailability:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Preferred pharmacy local'
        value: {
          qid: surveyDataset_SA:SA_RX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order Rx available'
        value: {
          qid: surveyDataset_SA:SA_RX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Other local pharmacy'
        value: {
          qid: surveyDataset_SA:SA_RX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx cost'
        value: {
          qid: surveyDataset_SA:SA_RX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Premium/Coverages Composite'
        value: {
          qid: PremiumCoverages:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand cost of plan (premium)'
        value: {
          qid: surveyDataset_SA:SA_PC1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand cost of care (deductable/copay/OOP max)'
        value: {
          qid: surveyDataset_SA:SA_PC2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Covered services'
        value: {
          qid: surveyDataset_SA:SA_PC3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Supplemental Benefits'
        value: {
          qid: surveyDataset_SA:SA_SB1
          target: 87
          removeEmptyRows: true
        }
      }
    }
    row cut #row {
      value: @selectorBackgroundVar1.selected
      showLabel: false
      total: "first"
      totalLabel: "Total"
    }
    removeEmptyRows: true

    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column #column_2 {
      cell microchart #cell {
        value: average(numeric(@selectorQuestion1.selected.qid))
        microchart bar #barMicrochart {
          valuePosition: outer
          colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          min: 0
          max: 100
        }
        format: OneDecimalNumberFormatter
        target: @selectorQuestion1.selected.target
      }
      label: "Score"
    }
    column #column_4 {
      cell #cell {
        value: @selectorQuestion1.selected.target
      }
      label: "PG Benchmark"
    }
    column #column_3 {
      cell #cell {
        value: average(numeric(@selectorQuestion1.selected.qid)) - @selectorQuestion1.selected.target
        format: OneDecimalNumberFormatter
      }
      label: "Gap to PG Benchmark"
    }
  }
  hide: false
  modal: true
}





page #SA_OA_Plus_Grid {
  widget dataGrid #dataGridWidget {
    cardCorners: '20px'
    label: "SALES KPI's"
    size: medium
    column cutByDate #column_2 {
      value: surveyDataset_SA:interview_end
      total: "none"
      showLabel: false
    }
    column cutByDate #column {
      label: " "
      value: surveyDataset_SA:interview_end
      showLabel: false
      total: "none"
      breakdownBy: "calendarMonth"
      align: true
      start: "-1 month"
    }
    row #row {
      cell #cell {
        value: average(numeric(surveyDataset_SA:OA1))
        showBase: true
        format: OneDecimalNumberFormatter
        view: comparativeStatisticView
      }
      label: "Overall Experience"
    }
    row #row_2 {
      cell #cell {
        value: average(numeric(ProviderAvailability:value))
        showBase: true
        view: comparativeStatisticView_2
        format: OneDecimalNumberFormatter
      }
      label: "Provider Availability"
    }
    row #row_3 {
      cell #cell {
        value: average(numeric(RxAvailability:value))
        showBase: false
        view: comparativeStatisticView_3
        format: OneDecimalNumberFormatter
      }
      label: "Rx Availability"
    }
    row #row_4 {
      cell #cell {
        value: average(numeric(PremiumCoverages:value))
        showBase: false
        view: comparativeStatisticView_4
        format: OneDecimalNumberFormatter
      }
      label: "Premium/Coverages"
    }
    row #row_5 {
      cell #cell {
        value: average(numeric(surveyDataset_SA:SA_SB1))
        showBase: false
        view: comparativeStatisticView_5
        format: OneDecimalNumberFormatter
      }
      label: "Supplemental benefits"
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    view comparativeStatistic #comparativeStatisticView_2 {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    view comparativeStatistic #comparativeStatisticView_3 {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    view comparativeStatistic #comparativeStatisticView_4 {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    view comparativeStatistic #comparativeStatisticView_5 {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    significanceTesting: true
    confidenceLevels: "95"
  }
  label: "SA_OA+ grid"
  hide: false
  modal: true
  modalSize: "medium"
}





page #SA_OA_trend_line {
  widget chart #SAtrendchart {
    cardCorners: '20px'
    label: "What are scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
        showBaseInTooltip: false
      }
      label: "Overall Experience with SALES"
      value: average(numeric(surveyDataset_SA:OA1))

      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Provider Availability"
      value: average(numeric(ProviderAvailability:value))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rx Availability"
      value: average(numeric(RxAvailability:value))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Premium/Coverages"
      value: average(numeric(PremiumCoverages:value))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Supplemental Benefits "
      value: average(numeric(surveyDataset_SA:SA_SB1))
      format: OneDecimalNumberFormatter
    }

    navigateTo: ""
    description: "SALES - Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "SA Composites trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_KDA_Correlation {
  label: "SA KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #MTM_SA_OA1_keyDriversWidget {
    cardCorners: '20px'
    label: "Sales Key Drivers of the Overall Experience Rating (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_SA:OA1
    independentVariables: surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8, surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4, surveyDataset_SA:SA_RX5, surveyDataset_SA:SA_RX6, surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3, surveyDataset_SA:SA_SB1
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 58
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    showModelDetails: true
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #FOUNDATIONS {





  label: "FOUNDATIONS"
  widget canvas #NP_KPI_scores_divider_canvasWidget {
    label: "NP KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "FOUNDATIONS KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #NP_KPI_scores_tabs_canvasWidget {
    label: "NP KPI scores tabs"
    container: container position {
      width: 1368px
      height: "58px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "845px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1183px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "6px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "7px"
        left: "1325px"
      }
      area #area_10 {
        position: "absolute"
        top: "33px"
        left: "309px"
      }
      area #area_12 {
        position: "absolute"
        top: "35px"
        left: "1170px"
      }
      area #area_13 {
        position: "absolute"
        top: "37px"
        left: "832px"
      }
    }
    tile text #MTM_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_NP.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    cardTransparent: true
    tile text #textTile {
      value: "Rating of Doctors"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Rating of Doctors"
      value: average(numeric(Doctors:value))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_NP:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_NPS_StackedBar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_DR_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_OA3_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_NP.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_NP.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_7 {
      areaId: "area_13"
      label: "Premium/Coverages"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_DR2) >= 0 OR numeric(surveyDataset_NP:NP_DR4) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #NPtrendchart_1 {
    cardCorners: '20px'
    label: "How is FOUNDATIONS NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_NP.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #NPtrendchart_3 {
    cardCorners: '20px'
    label: "How are FOUNDATIONS KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_NP:OA3))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Doctors"
      value: average(numeric(Doctors:value))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of PCP"
      value: average(numeric(surveyDataset_NP:NP_DR2))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Specialist"
      value: average(numeric(surveyDataset_NP:NP_DR4))
      format: OneDecimalNumberFormatter
    }


    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #NP_KDA_divider_canvasWidget {
    label: "NP Key Drivers of KPIs divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "FOUNDATIONS Key Drivers of KPIs"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget keyDrivers #NP_OA2_keyDriversWidget {
    cardCorners: '20px'
    label: "NPS"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_ACR1, surveyDataset_NP:NP_ACR2, surveyDataset_NP:NP_ACR3, surveyDataset_NP:NP_ACR4, surveyDataset_NP:NP_BC1, surveyDataset_NP:NP_BC2, surveyDataset_NP:NP_BC3, surveyDataset_NP:NP_PX1, surveyDataset_NP:NP_PX2, surveyDataset_NP:NP_PX3, surveyDataset_NP:NP_UP1, surveyDataset_NP:NP_UP2, surveyDataset_NP:NP_UP3, surveyDataset_NP:NP_UP4, surveyDataset_NP:NP_UP5, surveyDataset_NP:NP_UP6, surveyDataset_NP:NP_YH1, surveyDataset_NP:NP_YH2, surveyDataset_NP:NP_BI1, surveyDataset_NP:NP_BI2, surveyDataset_NP:NP_DR2, surveyDataset_NP:NP_DR4
  }
  widget keyDrivers #NP_OA3_keyDriversWidget {
    cardCorners: '20px'
    label: "Rating of Health Plan"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
    dependentVariable: surveyDataset_NP:OA3
    independentVariables: surveyDataset_NP:NP_ACR1, surveyDataset_NP:NP_ACR2, surveyDataset_NP:NP_ACR3, surveyDataset_NP:NP_ACR4, surveyDataset_NP:NP_BC1, surveyDataset_NP:NP_BC2, surveyDataset_NP:NP_BC3, surveyDataset_NP:NP_PX1, surveyDataset_NP:NP_PX2, surveyDataset_NP:NP_PX3, surveyDataset_NP:NP_UP1, surveyDataset_NP:NP_UP2, surveyDataset_NP:NP_UP3, surveyDataset_NP:NP_UP4, surveyDataset_NP:NP_UP5, surveyDataset_NP:NP_UP6, surveyDataset_NP:NP_YH1, surveyDataset_NP:NP_YH2, surveyDataset_NP:NP_BI1, surveyDataset_NP:NP_BI2, surveyDataset_NP:NP_DR2, surveyDataset_NP:NP_DR4
  }
  widget canvas #NP_SectionScores_divider_canvasWidget {
    label: "NP Section scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "FOUNDATIONS Section scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #NP_SectionTabs_canvasWidget {
    label: "NP Section scores tabs divider"
    container: container position {
      width: 1368px
      height: "57px"
      background: rgba(255, 255, 255, 0)
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "24px"
        left: "84px"
        position: "absolute"
      }
      area #area_9 {
        position: "absolute"
        top: "0px"
        left: "226px"
      }
      area #area_10 {
        position: "absolute"
        top: "24px"
        left: "310px"
      }
      area #area_11 {
        position: "absolute"
        top: "0px"
        left: "452px"
      }
      area #area_12 {
        position: "absolute"
        top: "24px"
        left: "536px"
      }
      area #area_13 {
        position: "absolute"
        top: "0px"
        left: "678px"
      }
      area #area_14 {
        position: "absolute"
        top: "24px"
        left: "762px"
      }
      area #area_15 {
        position: "absolute"
        top: "0px"
        left: "904px"
      }
      area #area_16 {
        position: "absolute"
        top: "24px"
        left: "988px"
      }
      area #area_17 {
        position: "absolute"
        top: "0px"
        left: "1131px"
      }
      area #area_18 {
        position: "absolute"
        top: "24px"
        left: "1215px"
      }
      area #area_19 {
        position: "absolute"
        top: "34px"
        left: "84px"
      }
      area #area_20 {
        position: "absolute"
        top: "35px"
        left: "310px"
      }
      area #area_21 {
        position: "absolute"
        top: "35px"
        left: "536px"
      }
      area #area_22 {
        position: "absolute"
        top: "35px"
        left: "762px"
      }
      area #area_23 {
        position: "absolute"
        top: "35px"
        left: "988px"
      }
      area #area_24 {
        position: "absolute"
        top: "35px"
        left: "1215px"
      }
      area #area_25 {
        position: "absolute"
        top: "6px"
        left: "184px"
      }
      area #area_26 {
        position: "absolute"
        top: "7px"
        left: "410px"
      }
      area #area_27 {
        position: "absolute"
        top: "7px"
        left: "635px"
      }
      area #area_28 {
        position: "absolute"
        top: "6px"
        left: "862px"
      }
      area #area_29 {
        position: "absolute"
        top: "6px"
        left: "1088px"
      }
      area #area_30 {
        position: "absolute"
        top: "7px"
        left: "1315px"
      }
    }
    cardTransparent: true

    tile text #NP_AC_textTile {
      value: "Access To Care"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "225px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Access To Care"
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "Access To Care"
      value: average(numeric(AccessToCare:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_5 {
      value: "Benefits and Coverage"
      areaId: "area_9"
      style #style {
        fontSize: 16
        width: "225px"
        height: "67px"
        textAlign: "left"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Benefits and Coverage"
    }
    tile value #valueTile_5 {
      areaId: "area_10"
      label: "Benefits and Coverage"
      value: average(numeric(BenefitsCoverage:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_6 {
      value: "Prescriptions"
      areaId: "area_11"
      style #style {
        fontSize: 16
        width: "225px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Prescriptions"
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "Prescriptions"
      value: average(numeric(Prescriptions:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_7 {
      value: "Using Your Health Plan"
      areaId: "area_13"
      style #style {
        fontSize: 16
        width: "225px"
        height: "67px"
        textAlign: "left"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Using Your Health Plan"
    }
    tile value #valueTile_7 {
      areaId: "area_14"
      label: "Using Your Health Plan"
      value: average(numeric(UsingHP:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_8 {
      value: "Your Health"
      areaId: "area_15"
      style #style {
        fontSize: 16
        width: "225px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Your Health"
    }
    tile value #valueTile_8 {
      areaId: "area_16"
      label: "Your Health"
      value: average(numeric(YourHealth:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_9 {
      value: "Brand Image"
      areaId: "area_17"
      style #style {
        fontSize: 16
        width: "225px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Brand Image"
    }
    tile value #valueTile_9 {
      areaId: "area_18"
      label: "Brand Image"
      value: average(numeric(BrandImage:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_10 {
      areaId: "area_19"
      label: "Access to Care"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_ACR1) >= 0 OR numeric(surveyDataset_NP:NP_ACR2) >= 0 OR numeric(surveyDataset_NP:NP_ACR3) >= 0 OR numeric(surveyDataset_NP:NP_ACR4) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_11 {
      areaId: "area_20"
      label: "Benefits and Coverages"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_BC1) >= 0 OR numeric(surveyDataset_NP:NP_BC2) >= 0 OR numeric(surveyDataset_NP:NP_BC3) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_12 {
      areaId: "area_21"
      label: "Prescriptions"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_PX1) >= 0 OR numeric(surveyDataset_NP:NP_PX2) >= 0 OR numeric(surveyDataset_NP:NP_PX3) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_13 {
      areaId: "area_22"
      label: "Using Your Health Plan"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_UP1) >= 0 OR numeric(surveyDataset_NP:NP_UP2) >= 0 OR numeric(surveyDataset_NP:NP_UP3) >= 0 OR numeric(surveyDataset_NP:NP_UP4) >= 0 OR numeric(surveyDataset_NP:NP_UP5) >= 0 OR numeric(surveyDataset_NP:NP_UP6) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_14 {
      areaId: "area_23"
      label: "Your Health"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_YH1) >= 0 OR numeric(surveyDataset_NP:NP_YH2) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_15 {
      areaId: "area_24"
      label: "Brand Image"
      value: count(surveyDataset_NP:respid, numeric(surveyDataset_NP:NP_BI1) >= 0 OR numeric(surveyDataset_NP:NP_BI2) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_25"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_AC_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_26"
      style #style {
        width: "34px"
        opacity: 1
      }
      navigateTo: "NP_BC_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_27"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_PX_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_28"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_UP_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_5 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_29"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_YH_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_6 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_30"
      style #style {
        width: "34px"
      }
      navigateTo: "NP_BI_stacked_bar"
      navigateOptions: "same_tab"
    }
  }
  widget chart #NPtrendchart_2 {
    cardCorners: '20px'
    label: "How are FOUNDATIONS Section scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Access to Care"
      value: average(numeric(AccessToCare:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Benefits and Coverage"
      value: average(numeric(BenefitsCoverage:value))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Prescriptions"
      value: average(numeric(Prescriptions:value))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Using Your Health Plan"
      value: average(numeric(UsingHP:value))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Your Health"
      value: average(numeric(YourHealth:value))
      format: OneDecimalNumberFormatter
    }
    series #series_6 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Brand Image"
      value: average(numeric(BrandImage:value))
      format: OneDecimalNumberFormatter
    }
    description: ""
    size: large
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #NP_ScoreComparison_divider {
    label: "NP Score Comparison Divider Canvas"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "5px"
        left: "63px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "FOUNDATIONS Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #NP_Top10_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_NP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_NP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_NP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_NP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_NP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_NP:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_NP:OA2
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_NP:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rating of Doctors Composite'
        value: {
          qid: Doctors:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rating of PCP'
        value: {
          qid: surveyDataset_NP:NP_DR2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rating of Specialist'
        value: {
          qid: surveyDataset_NP:NP_DR4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Access to Care Composite'
        value: {
          qid: AccessToCare:value
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of primary care doctors'
        value: {
          qid: surveyDataset_NP:NP_ACR1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of specialists'
        value: {
          qid: surveyDataset_NP:NP_ACR2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of labs/testing sites'
        value: {
          qid: surveyDataset_NP:NP_ACR3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of pharmacies'
        value: {
          qid: surveyDataset_NP:NP_ACR4
          target: 87
          removeEmptyRows: true
        }
      },      
      item {
        label: 'Benefits and Coverage Composite'
        value: {
          qid: BenefitsCoverage:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Coverage of doctor visits'
        value: {
          qid: surveyDataset_NP:NP_BC1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Coverage of labs/tests'
        value: {
          qid: surveyDataset_NP:NP_BC2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Value of benefits'
        value: {
          qid: surveyDataset_NP:NP_BC3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Prescriptions Composite'
        value: {
          qid: Prescriptions:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of obtaining Rx'
        value: {
          qid: surveyDataset_NP:NP_PX1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Cost of Rx'
        value: {
          qid: surveyDataset_NP:NP_PX2
          target: 87
          removeEmptyRows: true
        }
      },
            item {
        label: 'Coverage of Rx'
        value: {
          qid: surveyDataset_NP:NP_PX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Using Your Health Plan Composite'
        value: {
          qid: UsingHP:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of getting benefits info'
        value: {
          qid: surveyDataset_NP:NP_UP1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of getting provider info'
        value: {
          qid: surveyDataset_NP:NP_UP2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Wellness plan'
        value: {
          qid: surveyDataset_NP:NP_UP3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Plan rep response'
        value: {
          qid: surveyDataset_NP:NP_UP4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of sbumitting claim'
        value: {
          qid: surveyDataset_NP:NP_UP5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of reimbursement'
        value: {
          qid: surveyDataset_NP:NP_UP6
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Your Health Composite'
        value: {
          qid: YourHealth:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand your responsibilities in care'
        value: {
          qid: surveyDataset_NP:NP_YH1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Know what you can do to affect health'
        value: {
          qid: surveyDataset_NP:NP_YH2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Brand Image Composite'
        value: {
          qid: BrandImage:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Plan is market leader'
        value: {
          qid: surveyDataset_NP:NP_BI1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Plan is trustworthy'
        value: {
          qid: surveyDataset_NP:NP_BI2
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget chart #NP_Bottom10_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_NP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_NP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_NP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_NP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_NP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_NP:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_NP:OA2
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_NP:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rating of Doctors Composite'
        value: {
          qid: Doctors:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rating of PCP'
        value: {
          qid: surveyDataset_NP:NP_DR2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rating of Specialist'
        value: {
          qid: surveyDataset_NP:NP_DR4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Access to Care Composite'
        value: {
          qid: AccessToCare:value
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of primary care doctors'
        value: {
          qid: surveyDataset_NP:NP_ACR1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of specialists'
        value: {
          qid: surveyDataset_NP:NP_ACR2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of labs/testing sites'
        value: {
          qid: surveyDataset_NP:NP_ACR3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Availability of pharmacies'
        value: {
          qid: surveyDataset_NP:NP_ACR4
          target: 87
          removeEmptyRows: true
        }
      },      
      item {
        label: 'Benefits and Coverage Composite'
        value: {
          qid: BenefitsCoverage:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Coverage of doctor visits'
        value: {
          qid: surveyDataset_NP:NP_BC1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Coverage of labs/tests'
        value: {
          qid: surveyDataset_NP:NP_BC2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Value of benefits'
        value: {
          qid: surveyDataset_NP:NP_BC3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Prescriptions Composite'
        value: {
          qid: Prescriptions:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of obtaining Rx'
        value: {
          qid: surveyDataset_NP:NP_PX1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Cost of Rx'
        value: {
          qid: surveyDataset_NP:NP_PX2
          target: 87
          removeEmptyRows: true
        }
      },
            item {
        label: 'Coverage of Rx'
        value: {
          qid: surveyDataset_NP:NP_PX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Using Your Health Plan Composite'
        value: {
          qid: UsingHP:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of getting benefits info'
        value: {
          qid: surveyDataset_NP:NP_UP1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of getting provider info'
        value: {
          qid: surveyDataset_NP:NP_UP2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Wellness plan'
        value: {
          qid: surveyDataset_NP:NP_UP3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Plan rep response'
        value: {
          qid: surveyDataset_NP:NP_UP4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of sbumitting claim'
        value: {
          qid: surveyDataset_NP:NP_UP5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of reimbursement'
        value: {
          qid: surveyDataset_NP:NP_UP6
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Your Health Composite'
        value: {
          qid: YourHealth:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand your responsibilities in care'
        value: {
          qid: surveyDataset_NP:NP_YH1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Know what you can do to affect health'
        value: {
          qid: surveyDataset_NP:NP_YH2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Brand Image Composite'
        value: {
          qid: BrandImage:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Plan is market leader'
        value: {
          qid: surveyDataset_NP:NP_BI1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Plan is trustworthy'
        value: {
          qid: surveyDataset_NP:NP_BI2
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #NP_SectionComponent_divider {
    label: "NP Section and Component score Divider Canvas"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "5px"
        left: "60px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "FOUNDATIONS Section and Component Scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget headline #NP_AC_Dial {
    cardCorners: '20px'
    label: "Access to Care"
    tile gauge #gaugeTile {
      value: average(numeric(AccessToCare:value))
      format: OneDecimalNumberFormatter
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      targetFormat: OneDecimalNumberFormatter
      label: "Section Score"
      min: 0
      max: 100
      showRange: true
      navigateTo: "NP_AC_Components_stacked_bar"
      navigateOptions: "same_tab"
      target: 77
      belowTargetLabel: "Gap to PG Benchmark"
      aboveTargetLabel: "Avove PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_1__row {
        value: surveyDataset_NP:Dial__gridTile_1__variable$field
      }
      cell #Dial__gridTile_1__column__cell {
        value: average(numeric(surveyDataset_NP:Dial__gridTile_1__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_1__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_1__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: "auto"
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_1__column {
        hide: false
      }
      sort rows #Dial__gridTile_1__sort {
        sortBy: "/Dial__gridTile_1__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_1__row
        column: @Dial__gridTile_1__column
        cell: @Dial__gridTile_1__column__cell
        sort: @Dial__gridTile_1__sort
        variable: @Dial__gridTile_1__variable
        chartColumn: @Dial__gridTile_1__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "NP_AC_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "NP_AC_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "NP_AC_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Comment%20button.png"
      padding: true
      navigateTo: "NP_AC_Comments"
      navigateOptions: "same_tab"
    }
  }
  widget headline #NP_BC_Dial {
    cardCorners: '20px'
    label: "Benefits and Coverage"
    tile gauge #gaugeTile {
      value: average(numeric(BenefitsCoverage:value))
      format: OneDecimalNumberFormatter
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      targetFormat: OneDecimalNumberFormatter
      label: "Section Score"
      min: 0
      max: 100
      showRange: true
      navigateTo: "NP_BC_Components_stacked_bar"
      navigateOptions: "same_tab"
      target: 77
      belowTargetLabel: "Gap to PG Benchmark"
      aboveTargetLabel: "Avove PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_2__row {
        value: surveyDataset_NP:Dial__gridTile_2__variable$field
      }
      cell #Dial__gridTile_2__column__cell {
        value: average(numeric(surveyDataset_NP:Dial__gridTile_2__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_2__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_2__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: "auto"
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_2__column {
        hide: false
      }
      sort rows #Dial__gridTile_2__sort {
        sortBy: "/Dial__gridTile_2__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_2__row
        column: @Dial__gridTile_2__column
        cell: @Dial__gridTile_2__column__cell
        sort: @Dial__gridTile_2__sort
        variable: @Dial__gridTile_2__variable
        chartColumn: @Dial__gridTile_2__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "NP_BC_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "NP_BC_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "NP_BC_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Comment%20button.png"
      padding: true
      navigateTo: "NP_BC_Comments"
      navigateOptions: "same_tab"
    }
  }
  widget headline #NP_RX_Dial {
    cardCorners: '20px'
    label: "Prescriptions"
    tile gauge #gaugeTile {
      value: average(numeric(Prescriptions:value))
      format: OneDecimalNumberFormatter
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      targetFormat: OneDecimalNumberFormatter
      label: "Section Score"
      min: 0
      max: 100
      showRange: true
      navigateTo: "NP_PX_Components_stacked_bar"
      navigateOptions: "same_tab"
      target: 77
      belowTargetLabel: "Gap to PG Benchmark"
      aboveTargetLabel: "Avove PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_3__row {
        value: surveyDataset_NP:Dial__gridTile_3__variable$field
      }
      cell #Dial__gridTile_3__column__cell {
        value: average(numeric(surveyDataset_NP:Dial__gridTile_3__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_3__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_3__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: "auto"
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_3__column {
        hide: false
      }
      sort rows #Dial__gridTile_3__sort {
        sortBy: "/Dial__gridTile_3__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_3__row
        column: @Dial__gridTile_3__column
        cell: @Dial__gridTile_3__column__cell
        sort: @Dial__gridTile_3__sort
        variable: @Dial__gridTile_3__variable
        chartColumn: @Dial__gridTile_3__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "NP_PX_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "NP_PX_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "NP_PX_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Comment%20button.png"
      padding: true
      navigateTo: "NP_PX_Comments"
      navigateOptions: "same_tab"
    }
  }
  widget headline #NP_UP_Dial {
    cardCorners: '20px'
    label: "Using Your Health Plan"
    tile gauge #gaugeTile {
      value: average(numeric(UsingHP:value))
      format: OneDecimalNumberFormatter
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      targetFormat: OneDecimalNumberFormatter
      label: "Section Score"
      min: 0
      max: 100
      showRange: true
      navigateTo: "NP_UP_Components_stacked_bar"
      navigateOptions: "same_tab"
      target: 77
      belowTargetLabel: "Gap to PG Benchmark"
      aboveTargetLabel: "Avove PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_4__row {
        value: surveyDataset_NP:Dial__gridTile_4__variable$field
      }
      cell #Dial__gridTile_4__column__cell {
        value: average(numeric(surveyDataset_NP:Dial__gridTile_4__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_4__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_4__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: "auto"
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_4__column {
        hide: false
      }
      sort rows #Dial__gridTile_4__sort {
        sortBy: "/Dial__gridTile_4__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_4__row
        column: @Dial__gridTile_4__column
        cell: @Dial__gridTile_4__column__cell
        sort: @Dial__gridTile_4__sort
        variable: @Dial__gridTile_4__variable
        chartColumn: @Dial__gridTile_4__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "NP_UP_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "NP_UP_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "NP_UP_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Comment%20button.png"
      padding: true
      navigateTo: "NP_UP_Comments"
      navigateOptions: "same_tab"
    }
  }
  widget headline #NP_YH_Dial {
    cardCorners: '20px'
    label: "Your Health"
    tile gauge #gaugeTile {
      value: average(numeric(YourHealth:value))
      format: OneDecimalNumberFormatter
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      targetFormat: OneDecimalNumberFormatter
      label: "Section Score"
      min: 0
      max: 100
      showRange: true
      navigateTo: "NP_YH_Components_stacked_bar"
      navigateOptions: "same_tab"
      target: 77
      belowTargetLabel: "Gap to PG Benchmark"
      aboveTargetLabel: "Avove PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_5__row {
        value: surveyDataset_NP:Dial__gridTile_5__variable$field
      }
      cell #Dial__gridTile_5__column__cell {
        value: average(numeric(surveyDataset_NP:Dial__gridTile_5__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_5__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_5__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: "auto"
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_5__column {
        hide: false
      }
      sort rows #Dial__gridTile_5__sort {
        sortBy: "/Dial__gridTile_5__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_5__row
        column: @Dial__gridTile_5__column
        cell: @Dial__gridTile_5__column__cell
        sort: @Dial__gridTile_5__sort
        variable: @Dial__gridTile_5__variable
        chartColumn: @Dial__gridTile_5__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "NP_YH_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "NP_YH_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "NP_YH_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Comment%20button.png"
      padding: true
      navigateTo: "NP_YH_Comments"
      navigateOptions: "same_tab"
    }
  }
  widget headline #NP_BI_Dial {
    cardCorners: '20px'
    label: "Brand Image"
    tile gauge #gaugeTile {
      value: average(numeric(BrandImage:value))
      format: OneDecimalNumberFormatter
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      targetFormat: OneDecimalNumberFormatter
      label: "Section Score"
      min: 0
      max: 100
      showRange: true
      navigateTo: "NP_BI_Components_stacked_bar"
      navigateOptions: "same_tab"
      target: 77
      belowTargetLabel: "Gap to PG Benchmark"
      aboveTargetLabel: "Avove PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_6__row {
        value: surveyDataset_NP:Dial__gridTile_6__variable$field
      }
      cell #Dial__gridTile_6__column__cell {
        value: average(numeric(surveyDataset_NP:Dial__gridTile_6__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_6__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_6__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: "auto"
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_6__column {
        hide: false
      }
      sort rows #Dial__gridTile_6__sort {
        sortBy: "/Dial__gridTile_6__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_6__row
        column: @Dial__gridTile_6__column
        cell: @Dial__gridTile_6__column__cell
        sort: @Dial__gridTile_6__sort
        variable: @Dial__gridTile_6__variable
        chartColumn: @Dial__gridTile_6__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "NP_BI_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "NP_BI_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "NP_BI_KDA_Correlation"
      navigateOptions: "same_tab"
    }
  }
  widget canvas #NP_Comment_divider {
    label: "NP Comments Divider Canvas"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "5px"
        left: "63px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall FOUNDATIONS experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #NP_Comments {
    cardCorners: '20px'
    label: "Please describe a good or bad experience"
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_NP:OA4 != ""
      }
      comment: surveyDataset_NP:OA4
    }
    size: large
    table: surveyDataset_NP:
    cardBackground: #ffffff
    column value #NP_OA3_valueColumn {
      label: "Rating of Health Plan Response"
      value: surveyDataset_NP.response:OA3
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Rating of Health Plan Score"
      value: average(numeric(surveyDataset_NP.response:OA3))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #NP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_NP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_NP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_NP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #NP_Response_divider {
    label: "NP Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "5px"
        left: "64px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "FOUNDATIONS Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #NP_surveyMetricsWidget {
    cardCorners: '20px'
    label: "FOUNDATIONS Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_NP
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1
}





page #NP_NPS_StackedBar {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "FOUNDATIONS NPS"
    series #series {
      value: count(surveyDataset_NP.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_NP:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "How likely is it that you would recommend your health plan to a friend or colleague?"
    layout: "vertical"
  }
  widget headline #NP_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_NP.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_NP.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #NP_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_NP.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_NP.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #NP_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_NP.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_NP.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "NP_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #NP_DR_stacked_bar {
  widget chart #NP_DR_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rating of Doctors"
    series #series {
      value: count(Doctors:value)
      label: "Dr. Rating"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: Doctors:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
  }
  widget chart #NP_DR_stacked_bar_COMPONENTS_chartWidget {
    cardCorners: '20px'
    label: "Rating of Doctors Components"
    series #series {
      value: count(Doctors:value)
      label: "Dr. Rating"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: Doctors:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    category cut #cutCategory {
      value: Doctors:field
    }
  }
  label: "NP_DRs stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #NP_OA3_stacked_bar {
  widget chart #NP_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "FOUNDATIONS - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_NP.response:OA3)
      label: "RHP"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_NP:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }

  label: "NP_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #NP_AC_stacked_bar {
  label: "NP_AC stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #NP_AC_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Access to Care"
    series #series {
      value: count(AccessToCare:value)
      label: "Access To Care"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: AccessToCare:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #NP_AC_Components_stacked_bar {
  label: "NP_AC Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #NP_AC_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Access to Care Components"
    series #series {
      value: count(AccessToCare:value)
      label: "Access to Care"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: AccessToCare:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: AccessToCare:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #NP_AC_grid {
  label: "NP_AC grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #NP_AC_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(AccessToCare:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_NP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: AccessToCare:field
      showLabel: false
      totalLabel: "Access to Care"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #NP_AC_trend_line {
  widget chart #NPtrendchart {
    cardCorners: '20px'
    label: "What are FOUNDATIONS - Access to Care scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Access to Care"
      value: average(numeric(AccessToCare:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Availability of primary care doctors"
      value: average(numeric(surveyDataset_NP:NP_ACR1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Availability of specialists"
      value: average(numeric(surveyDataset_NP:NP_ACR2))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Availability of labs/testing sites"
      value: average(numeric(surveyDataset_NP:NP_ACR3))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Availability of pharmacies"
      value: average(numeric(surveyDataset_NP:NP_ACR4))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "FOUNDATIONS - AC Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "NP_AC trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_AC_KDA_Correlation {
  label: "NP_AC KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #NP_OA2_AC_keyDriversWidget {
    cardCorners: '20px'
    label: "Access to Care Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.61
    importanceLimit: -0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_ACR1, surveyDataset_NP:NP_ACR2, surveyDataset_NP:NP_ACR3, surveyDataset_NP:NP_ACR4
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #NP_AC_Comments {
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please describe a good or bad Access to Care experience "
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_NP:NP_AC5 != ""
      }
      comment: surveyDataset_NP:NP_AC5
    }
    size: large
    table: surveyDataset_NP:
    cardBackground: #ffffff
    column value #NP_AC1_valueColumn {
      label: "Availability of PCPs Response"
      value: surveyDataset_NP.response:NP_ACR1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_AC2_valueColumn {
      label: "Availability of Specialists Response"
      value: surveyDataset_NP.response:NP_ACR2
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_AC3_valueColumn {
      label: "Availability of labs/testing sites Response"
      value: surveyDataset_NP.response:NP_ACR3
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_AC4_valueColumn {
      label: "Availability of Pharmacies Response"
      value: surveyDataset_NP.response:NP_ACR4
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_NP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_NP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_NP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  label: "NP_AC Comments"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_BC_stacked_bar {
  label: "NP_BC stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #NP_BC_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Benefits and Coverage"
    series #series {
      value: count(BenefitsCoverage:value)
      label: "Benefits and Coverage"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: BenefitsCoverage:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #NP_BC_Components_stacked_bar {
  label: "NP_BC Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #NP_BC_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Benefits and Coverage Components"
    series #series {
      value: count(BenefitsCoverage:value)
      label: "Benefits and Coverage"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: BenefitsCoverage:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: BenefitsCoverage:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #NP_BC_grid {
  label: "NP_BC grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #NP_BC_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(BenefitsCoverage:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_NP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: BenefitsCoverage:field
      showLabel: false
      totalLabel: "Benefits and Coverage"
      label: " "
    }

    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #NP_BC_trend_line {
  widget chart #NPtrendchart {
    cardCorners: '20px'
    label: "What are FOUNDATIONS - Benefits and Coverage scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Benefits and Coverage"
      value: average(numeric(BenefitsCoverage:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Coverage of doctor visits"
      value: average(numeric(surveyDataset_NP:NP_BC1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Coverage of labs/tests"
      value: average(numeric(surveyDataset_NP:NP_BC2))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Value of benefits"
      value: average(numeric(surveyDataset_NP:NP_BC3))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "FOUNDATIONS - BC Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "NP_BC trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_BC_KDA_Correlation {
  label: "NP_BC KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #NP_OA2_BC_keyDriversWidget {
    cardCorners: '20px'
    label: "Benefits and Coverage Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.57
    importanceLimit: 0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_BC1, surveyDataset_NP:NP_BC2, surveyDataset_NP:NP_BC3
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #NP_BC_Comments {
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please describe a good or bad Benefits and Coverage experience "
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_NP:NP_BC4 != ""
      }
      comment: surveyDataset_NP:NP_BC4
    }
    size: large
    table: surveyDataset_NP:
    cardBackground: #ffffff
    column value #NP_BC1_valueColumn {
      label: "Coverage of doctor visits Response"
      value: surveyDataset_NP.response:NP_BC1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_BC2_valueColumn {
      label: "Coverage of labs/tests Response"
      value: surveyDataset_NP.response:NP_BC2
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_BC3_valueColumn {
      label: "Value of benefits Response"
      value: surveyDataset_NP.response:NP_BC3
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_NP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_NP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_NP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  label: "NP_BC Comments"
  hide: false
  modal: true
  modalSize: "large"
}




page #NP_PX_stacked_bar {
  label: "NP_PX stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #NP_PX_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Prescriptions"
    series #series {
      value: count(Prescriptions:value)
      label: "Prescriptions"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: Prescriptions:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #NP_PX_Components_stacked_bar {
  label: "NP_PX Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #NP_PX_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Prescriptions Components"
    series #series {
      value: count(Prescriptions:value)
      label: "Prescriptions"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: Prescriptions:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: Prescriptions:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #NP_PX_grid {
  label: "NP_PX grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #NP_PX_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(Prescriptions:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_NP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: Prescriptions:field
      showLabel: false
      totalLabel: "Prescriptions"
      label: " "
    }

    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #NP_PX_trend_line {
  widget chart #NPtrendchart {
    cardCorners: '20px'
    label: "What are FOUNDATIONS - Prescriptions scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Prescriptions"
      value: average(numeric(Prescriptions:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Ease of obtaining prescriptions"
      value: average(numeric(surveyDataset_NP:NP_PX1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Cost of prescriptions"
      value: average(numeric(surveyDataset_NP:NP_PX2))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Coverage of prescribed medications"
      value: average(numeric(surveyDataset_NP:NP_PX3))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "FOUNDATIONS - PX Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "NP_PX trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_PX_KDA_Correlation {
  label: "NP_PX KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #NP_OA2_PX_keyDriversWidget {
    cardCorners: '20px'
    label: "Prescriptions Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.33
    importanceLimit: 0.04
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_PX1, surveyDataset_NP:NP_PX2, surveyDataset_NP:NP_PX3
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #NP_PX_Comments {
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please describe a good or bad Prescriptions experience "
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_NP:NP_PX4 != ""
      }
      comment: surveyDataset_NP:NP_PX4
    }
    size: large
    table: surveyDataset_NP:
    cardBackground: #ffffff
    column value #NP_PX1_valueColumn {
      label: "Ease of obtaing prescriptions Response"
      value: surveyDataset_NP.response:NP_PX1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PX2_valueColumn {
      label: "Cost of prescriptions Response"
      value: surveyDataset_NP.response:NP_PX2
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PX3_valueColumn {
      label: "Coverage of prescribed medications Response"
      value: surveyDataset_NP.response:NP_PX3
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_NP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_NP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_NP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  label: "NP_PX Comments"
  hide: false
  modal: true
  modalSize: "large"
}




page #NP_UP_stacked_bar {
  label: "NP_UP stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #NP_UP_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Using Your Health Plan"
    series #series {
      value: count(UsingHP:value)
      label: "Using Your Health Plan"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: UsingHP:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #NP_UP_Components_stacked_bar {
  label: "NP_UP Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #NP_UP_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Using Your Health Plan Components"
    series #series {
      value: count(UsingHP:value)
      label: "Using Your Health Plan"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: UsingHP:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: UsingHP:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #NP_UP_grid {
  label: "NP_UP grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #NP_UP_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(UsingHP:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_NP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: UsingHP:field
      showLabel: false
      totalLabel: "Using Your Health Plan"
      label: " "
    }

    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #NP_UP_trend_line {
  widget chart #NPtrendchart {
    cardCorners: '20px'
    label: "What are FOUNDATIONS - Using Your Health Plan scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Using Your Health Plan"
      value: average(numeric(UsingHP:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Ease of getting benefits information"
      value: average(numeric(surveyDataset_NP:NP_UP1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Ease of getting provider information"
      value: average(numeric(surveyDataset_NP:NP_UP2))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Wellness plan"
      value: average(numeric(surveyDataset_NP:NP_UP3))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Plan rep's response to questions"
      value: average(numeric(surveyDataset_NP:NP_UP4))
      format: OneDecimalNumberFormatter
    }
    series #series_6 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Ease of submitting a claim"
      value: average(numeric(surveyDataset_NP:NP_UP5))
      format: OneDecimalNumberFormatter
    }
    series #series_7 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Timeliness of reimbursement"
      value: average(numeric(surveyDataset_NP:NP_UP6))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "FOUNDATIONS - UP Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "NP_UP trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_UP_KDA_Correlation {
  label: "NP_UP KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #NP_OA2_UP_keyDriversWidget {
    cardCorners: '20px'
    label: "Using Your Health Plan Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 51.28
    importanceLimit: 0.02
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_UP1, surveyDataset_NP:NP_UP2, surveyDataset_NP:NP_UP3, surveyDataset_NP:NP_UP4, surveyDataset_NP:NP_UP5, surveyDataset_NP:NP_UP6
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #NP_UP_Comments {
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please describe a good or bad Using Your Health Plan experience "
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_NP:NP_UP7 != ""
      }
      comment: surveyDataset_NP:NP_UP7
    }
    size: large
    table: surveyDataset_NP:
    cardBackground: #ffffff
    column value #NP_UP1_valueColumn {
      label: "Ease of getting benefits information Response"
      value: surveyDataset_NP.response:NP_UP1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_UP2_valueColumn {
      label: "Ease of getting provider information Response"
      value: surveyDataset_NP.response:NP_UP2
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_UP3_valueColumn {
      label: "Wellness plan Response"
      value: surveyDataset_NP.response:NP_UP3
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_UP4_valueColumn {
      label: "Plan rep's response to questions Response"
      value: surveyDataset_NP.response:NP_UP4
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_UP5_valueColumn {
      label: "Ease of submitting a claim Response"
      value: surveyDataset_NP.response:NP_UP5
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_UP6_valueColumn {
      label: "Timeliness of reimbursement Response"
      value: surveyDataset_NP.response:NP_UP6
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_NP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_NP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_NP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  label: "NP_UP Comments"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_YH_stacked_bar {
  label: "NP_YH stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #NP_YH_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Your Health"
    series #series {
      value: count(YourHealth:value)
      label: "Your Health"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: YourHealth:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #NP_YH_Components_stacked_bar {
  label: "NP_YH Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #NP_YH_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Your Health Components"
    series #series {
      value: count(YourHealth:value)
      label: "Your Health"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: YourHealth:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: YourHealth:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #NP_YH_grid {
  label: "NP_YH grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #NP_YH_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(YourHealth:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_NP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: YourHealth:field
      showLabel: false
      totalLabel: "Your Health"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #NP_YH_trend_line {
  widget chart #NPtrendchart {
    cardCorners: '20px'
    label: "What are FOUNDATIONS - Your Health scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Your Health"
      value: average(numeric(YourHealth:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Understand your responsibilities in care"
      value: average(numeric(surveyDataset_NP:NP_YH1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Know what you can do to affect your health"
      value: average(numeric(surveyDataset_NP:NP_YH2))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "FOUNDATIONS - YH Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "NP_YH trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_YH_KDA_Correlation {
  label: "NP_YH KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #NP_OA2_YH_keyDriversWidget {
    cardCorners: '20px'
    label: "Your Health Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.5
    importanceLimit: -0.02
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_YH1, surveyDataset_NP:NP_YH2
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #NP_YH_Comments {
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please describe a good or bad Your Health experience "
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_NP:NP_YH3 != ""
      }
      comment: surveyDataset_NP:NP_YH3
    }
    size: large
    table: surveyDataset_NP:
    cardBackground: #ffffff
    column value #NP_YH1_valueColumn {
      label: "Understand your responsibilities in care Response"
      value: surveyDataset_NP.response:NP_YH1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_YH2_valueColumn {
      label: "Know what you can do to affect your health Response"
      value: surveyDataset_NP.response:NP_YH2
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_NP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_NP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #NP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_NP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  label: "NP_YH Comments"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_BI_stacked_bar {
  label: "NP_BI stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #NP_BI_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Brand Image"
    series #series {
      value: count(BrandImage:value)
      label: "Brand Image"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: BrandImage:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #NP_BI_Components_stacked_bar {
  label: "NP_BI Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #NP_BI_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Brand Image Components"
    series #series {
      value: count(BrandImage:value)
      label: "Brand Image"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: BrandImage:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: BrandImage:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #NP_BI_grid {
  label: "NP_BI grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #NP_BI_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(BrandImage:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_NP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: BrandImage:field
      showLabel: false
      totalLabel: "Brand Image"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #NP_BI_trend_line {
  widget chart #NPtrendchart {
    cardCorners: '20px'
    label: "What are FOUNDATIONS - Brand Image scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Brand Image"
      value: average(numeric(BrandImage:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_NP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Health Plan is a market leader"
      value: average(numeric(surveyDataset_NP:NP_BI1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Health Plan is trustworthy"
      value: average(numeric(surveyDataset_NP:NP_BI2))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "FOUNDATIONS - BI Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "NP_BI trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #NP_BI_KDA_Correlation {
  label: "NP_BI KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #NP_OA2_BI_keyDriversWidget {
    cardCorners: '20px'
    label: "Brand Image Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.55
    importanceLimit: -0.07
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    dependentVariable: surveyDataset_NP:OA2
    independentVariables: surveyDataset_NP:NP_BI1, surveyDataset_NP:NP_BI2
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}






page #SALES {





  label: "SALES"
  widget canvas #SA_KPI_scores_divider {
    label: "SA KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #SA_KPIScores_tabs_divider {
    label: "SA KPI scores tabs divider"
    container: container position {
      width: 1368px
      height: "55px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "845px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1183px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "7px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "6px"
        left: "1326px"
      }
      area #area_10 {
        top: "32px"
        left: "309px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "832px"
      }
      area #area_12 {
        position: "absolute"
        top: "34px"
        left: "1170px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Overall Experience"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #SA_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_SA.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: average(numeric(surveyDataset_SA:OA1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_SA:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_OA2_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_OA1_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_OA3_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_SA.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_SA.response:OA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_SA.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #SA_NPS_trendchart {
    cardCorners: '20px'
    label: "How is SALES NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_SA.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #SA_KPI_trendchart {
    cardCorners: '20px'
    label: "How are SALES KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Overall Experience with SALES"
      value: average(numeric(surveyDataset_SA:OA1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_SA:OA3))
      format: OneDecimalNumberFormatter
    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #SA_KeyDrivers_divider {
    label: "SA Key Drivers of KPIs divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Key Drivers of KPIs"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget keyDrivers #SA_OA2_keyDriversWidget {
    cardCorners: '20px'
    label: "NPS"
    size: medium
    dependentVariable: surveyDataset_SA:OA2
    independentVariables: surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8, surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX6, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4, surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3, surveyDataset_SA:SA_SB1
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 48.48
    importanceLimit: 0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #SA_OA1_keyDriversWidget {
    cardCorners: '20px'
    label: "Overall Experience"
    size: small
    dependentVariable: surveyDataset_SA:OA1
    independentVariables: surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8, surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX6, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4, surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3, surveyDataset_SA:SA_SB1
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 48.48
    importanceLimit: 0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #SA_OA3_keyDriversWidget {
    cardCorners: '20px'
    label: "Rating of Health Plan"
    size: small
    dependentVariable: surveyDataset_SA:OA3
    independentVariables: surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8, surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX6, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4, surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3, surveyDataset_SA:SA_SB1
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 48.48
    importanceLimit: 0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget canvas #SA_Section_scores_divider {
    label: "SA Section scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Section scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #SA_SectionScores_tabs_divider {
    label: "SA Section scores tabs divider"
    container: container position {
      width: 1368px
      height: "59px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "687px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "140px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "17px"
        left: "840px"
        position: "absolute"
      }
      area #area_6 {
        top: "17px"
        left: "1183px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "0px"
        left: "343px"
      }
      area #area_8 {
        top: "22px"
        left: "483px"
        position: "absolute"
      }
      area #area_9 {
        position: "absolute"
        top: "35px"
        left: "140px"
      }
      area #area_10 {
        position: "absolute"
        top: "34px"
        left: "483px"
      }
      area #area_11 {
        position: "absolute"
        top: "35px"
        left: "827px"
      }
      area #area_12 {
        position: "absolute"
        top: "35px"
        left: "1170px"
      }
      area #area_13 {
        position: "absolute"
        top: "6px"
        left: "297px"
      }
      area #area_14 {
        position: "absolute"
        top: "7px"
        left: "639px"
      }
      area #area_15 {
        position: "absolute"
        top: "7px"
        left: "984px"
      }
      area #area_16 {
        position: "absolute"
        top: "8px"
        left: "1328px"
      }
    }
    cardTransparent: true

    tile text #SA_PA_textTile {
      value: "Provider Availability"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Provider Availability"
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "Provider Availability"
      value: average(numeric(ProviderAvailability:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_9"
      label: "Provider Availability"
      value: count(surveyDataset_SA:respid, numeric(surveyDataset_SA:SA_PA2) >= 0 OR numeric(surveyDataset_SA:SA_PA4) >= 0 OR numeric(surveyDataset_SA:SA_PA5) >= 0 OR numeric(surveyDataset_SA:SA_PA6) >= 0 OR numeric(surveyDataset_SA:SA_PA7) >= 0 OR numeric(surveyDataset_SA:SA_PA8) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_4 {
      value: "Rx Availability"
      areaId: "area_7"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Rx Availability"
    }
    tile value #valueTile_4 {
      areaId: "area_8"
      label: "Rx Availability"
      value: average(numeric(RxAvailability:value))
      style #style {
        fontSize: 16
        fontWeight: "bold"
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
      }
      valueFormatter: OneDecimalNumberFormatter
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      view: valueDefaultView
      formatString: "{value}"
    }

    tile value #valueTile_6 {
      areaId: "area_10"
      label: "Rx Availability"
      value: count(surveyDataset_SA:respid, numeric(surveyDataset_SA:SA_RX2) >= 0 OR numeric(surveyDataset_SA:SA_RX3) >= 0 OR numeric(surveyDataset_SA:SA_RX4) >= 0 OR numeric(surveyDataset_SA:SA_RX5) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile {
      value: "Premium/Coverages"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Premium/Coverages"
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Premium/Coverages"
      value: average(numeric(PremiumCoverages:value))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_7 {
      areaId: "area_11"
      label: "Premium/Coverages"
      value: count(surveyDataset_SA:respid, numeric(surveyDataset_SA:SA_PC1) >= 0 OR numeric(surveyDataset_SA:SA_PC2) >= 0 OR numeric(surveyDataset_SA:SA_PC3) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_3 {
      value: "Supplemental Benefits"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Supplemental Benefits"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "Supplemental Benefits"
      value: average(numeric(surveyDataset_SA:SA_SB1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_8 {
      areaId: "area_12"
      label: "Supplemental Benefits"
      value: count(surveyDataset_SA:respid, numeric(surveyDataset_SA:SA_SB1) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_13"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_PA_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_14"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_RX_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_15"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_PC_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_16"
      style #style {
        width: "34px"
      }
      navigateTo: "SA_SB1_stacked_bar"
      navigateOptions: "same_tab"
    }
  }
  widget chart #SA_SectionScore_trendchart {
    cardCorners: '20px'
    label: "How are SALES Section scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Provider Availability"
      value: average(numeric(ProviderAvailability:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rx Availability"
      value: average(numeric(RxAvailability:value))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Premium/Coverages"
      value: average(numeric(PremiumCoverages:value))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Supplemental Benefits "
      value: average(numeric(surveyDataset_SA:SA_SB1))
      format: OneDecimalNumberFormatter
    }


    description: ""
    size: large
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #SA_ScoreComparison_divider {
    label: "SA Score Comparison divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_SA:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_SA:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_SA:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_SA:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_SA:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_SA:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_SA:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_SA.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_SA:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Provider Availability Composite'
        value: {
          qid: ProviderAvailability:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Existing PCP in network'
        value: {
          qid: surveyDataset_SA:SA_PA2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Existing spec in network'
        value: {
          qid: surveyDataset_SA:SA_PA4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Hospital/facility in network'
        value: {
          qid: surveyDataset_SA:SA_PA5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'PCP local'
        value: {
          qid: surveyDataset_SA:SA_PA6
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Spec local'
        value: {
          qid: surveyDataset_SA:SA_PA7
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Finding provider(s) that meet certain characteristics'
        value: {
          qid: surveyDataset_SA:SA_PA8
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Pharmacy/Rx Availability Composite'
        value: {
          qid: RxAvailability:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Preferred pharmacy local'
        value: {
          qid: surveyDataset_SA:SA_RX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order Rx available'
        value: {
          qid: surveyDataset_SA:SA_RX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Other local pharmacy'
        value: {
          qid: surveyDataset_SA:SA_RX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx cost'
        value: {
          qid: surveyDataset_SA:SA_RX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Premium/Coverages Composite'
        value: {
          qid: PremiumCoverages:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand cost of plan (premium)'
        value: {
          qid: surveyDataset_SA:SA_PC1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand cost of care (deductable/copay/OOP max)'
        value: {
          qid: surveyDataset_SA:SA_PC2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Covered services'
        value: {
          qid: surveyDataset_SA:SA_PC3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Supplemental Benefits'
        value: {
          qid: surveyDataset_SA:SA_SB1
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: false
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget chart #SA_ScoreComparison_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_SA:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_SA:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_SA:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_SA:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_SA:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_SA:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_SA:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
      item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_SA.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
      item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_SA:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Provider Availability Composite'
        value: {
          qid: ProviderAvailability:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Existing PCP in network'
        value: {
          qid: surveyDataset_SA:SA_PA2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Existing spec in network'
        value: {
          qid: surveyDataset_SA:SA_PA4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Hospital/facility in network'
        value: {
          qid: surveyDataset_SA:SA_PA5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'PCP local'
        value: {
          qid: surveyDataset_SA:SA_PA6
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Spec local'
        value: {
          qid: surveyDataset_SA:SA_PA7
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Finding provider(s) that meet certain characteristics'
        value: {
          qid: surveyDataset_SA:SA_PA8
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Pharmacy/Rx Availability Composite'
        value: {
          qid: RxAvailability:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Preferred pharmacy local'
        value: {
          qid: surveyDataset_SA:SA_RX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order Rx available'
        value: {
          qid: surveyDataset_SA:SA_RX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Other local pharmacy'
        value: {
          qid: surveyDataset_SA:SA_RX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx cost'
        value: {
          qid: surveyDataset_SA:SA_RX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Premium/Coverages Composite'
        value: {
          qid: PremiumCoverages:value
          target: 55
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand cost of plan (premium)'
        value: {
          qid: surveyDataset_SA:SA_PC1
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Understand cost of care (deductable/copay/OOP max)'
        value: {
          qid: surveyDataset_SA:SA_PC2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Covered services'
        value: {
          qid: surveyDataset_SA:SA_PC3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Supplemental Benefits'
        value: {
          qid: surveyDataset_SA:SA_SB1
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #SA_SectionCompoenentScores_divider {
    label: "SA Section and Component Scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Section and Component Scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget headline #SA_PA_Dial {
    cardCorners: '20px'
    label: "Provider Availability"
    tile gauge #gaugeTile {
      value: average(numeric(ProviderAvailability:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "SA_PA_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"

    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_8__row {
        value: surveyDataset_SA:Dial__gridTile_8__variable$field

      }
      cell #Dial__gridTile_8__column__cell {
        value: average(numeric(surveyDataset_SA:Dial__gridTile_8__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_8__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_8__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_8__column {
        hide: false
      }
      sort rows #Dial__gridTile_8__sort {
        sortBy: "/Dial__gridTile_8__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_8__row
        column: @Dial__gridTile_8__column
        cell: @Dial__gridTile_8__column__cell
        sort: @Dial__gridTile_8__sort
        variable: @Dial__gridTile_8__variable
        chartColumn: @Dial__gridTile_8__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "SA_PA_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "SA_PA_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "SA_PA_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button.png"
      padding: true
      navigateTo: "SA_PA_Drilldown"
      navigateOptions: "same_tab"
    }
  }
  widget headline #SA_RX_Dial {
    cardCorners: '20px'
    label: "Rx Availability"
    tile gauge #gaugeTile {
      value: average(numeric(RxAvailability:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "SA_RX_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_9__row {

        value: surveyDataset_SA:Dial__gridTile_9__variable$field
      }
      cell #Dial__gridTile_9__column__cell {
        format: OneDecimalNumberFormatter
        value: average(numeric(surveyDataset_SA:Dial__gridTile_9__variable$value))
      }
      column #Dial__gridTile_9__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_9__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_9__column {
        hide: false
      }
      sort rows #Dial__gridTile_9__sort {
        sortBy: "/Dial__gridTile_9__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_9__row
        column: @Dial__gridTile_9__column
        cell: @Dial__gridTile_9__column__cell
        sort: @Dial__gridTile_9__sort
        variable: @Dial__gridTile_9__variable
        chartColumn: @Dial__gridTile_9__chartColumn
      }

    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      navigateTo: "SA_RX_grid"
      navigateOptions: "same_tab"
      padding: true
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      navigateTo: "SA_RX_trend_line"
      navigateOptions: "same_tab"
      padding: true
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "SA_RX_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button.png"
      padding: true
      navigateTo: "SA_RX_Drilldown"
      navigateOptions: "same_tab"
    }
  }
  widget headline #SA_PC_Dial {
    cardCorners: '20px'
    label: "Premium/Coverages"
    tile gauge #gaugeTile {
      value: average(numeric(PremiumCoverages:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "SA_PC_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_10__row {

        value: surveyDataset_SA:Dial__gridTile_10__variable$field
      }
      cell #Dial__gridTile_10__column__cell {
        format: OneDecimalNumberFormatter
        value: average(numeric(surveyDataset_SA:Dial__gridTile_10__variable$value))
      }
      column #Dial__gridTile_10__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_10__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_10__column {
        hide: false
      }
      sort rows #Dial__gridTile_10__sort {
        sortBy: "/Dial__gridTile_10__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_10__row
        column: @Dial__gridTile_10__column
        cell: @Dial__gridTile_10__column__cell
        sort: @Dial__gridTile_10__sort
        variable: @Dial__gridTile_10__variable
        chartColumn: @Dial__gridTile_10__chartColumn
      }

    }
    size: small
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      navigateTo: "SA_PC_grid"
      navigateOptions: "same_tab"
      padding: true
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "SA_PC_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      navigateTo: "SA_PC_SB_KDA_Correlation"
      navigateOptions: "same_tab"
      padding: true
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button.png"
      navigateTo: "SA_PC_Drilldown"
      navigateOptions: "same_tab"
      padding: true
    }
  }
  widget headline #SA_SB1_Dial {
    cardCorners: '20px'
    label: "Supplemental Benefits"
    tile gauge #gaugeTile {
      value: average(numeric(surveyDataset_SA:SA_SB1))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "SA_SB1_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"
    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_11__row {

        value: surveyDataset_SA:Dial__gridTile_11__variable$field
      }
      cell #Dial__gridTile_11__column__cell {
        format: OneDecimalNumberFormatter
        value: average(numeric(surveyDataset_SA:Dial__gridTile_11__variable$value))
      }
      column #Dial__gridTile_11__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_11__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_11__column {
        hide: false
      }
      sort rows #Dial__gridTile_11__sort {
        sortBy: "/Dial__gridTile_11__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_11__row
        column: @Dial__gridTile_11__column
        cell: @Dial__gridTile_11__column__cell
        sort: @Dial__gridTile_11__sort
        variable: @Dial__gridTile_11__variable
        chartColumn: @Dial__gridTile_11__chartColumn
      }
    }
    size: small
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      navigateTo: "SA_SB_grid"
      navigateOptions: "same_tab"
      padding: true
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "SA_SB_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      navigateTo: "SA_PC_SB_KDA_Correlation"
      navigateOptions: "same_tab"
      padding: true
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button.png"
      navigateTo: "SA_SB_Drilldown"
      navigateOptions: "same_tab"
      padding: true
    }
  }
  widget canvas #SA_Comment_divider {
    label: "SA Comment divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall SALES experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please provide any additional comments."
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_SA:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:OA4 != ""
      }
      comment: surveyDataset_SA:OA4
    }
    size: large
    table: surveyDataset_SA:
    cardBackground: #ffffff
    column value #SA_OA1_valueColumn {
      label: "Overall Experience Response"
      value: surveyDataset_SA.response:OA1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_SA.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #SA_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_SA.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #SA_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_SA.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #SA_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_SA.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #SA_Response_divider {
    label: "SA Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #SA_surveyMetricsWidget {
    cardCorners: '20px'
    label: "SALES Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_SA
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_OA1, fromQuestionFilter_CX_MEMST
}





page #SA_OA2_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "SALES NPS"
    series #series {
      value: count(surveyDataset_SA.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "On a scale of 0 to 10, how likely are you to recommend this health plan to a friend or a colleague?"
    layout: "vertical"
  }
  widget headline #SA_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_SA.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_SA.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #SA_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_SA.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_SA.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #SA_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_SA.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_SA.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "SA_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #SA_OA1_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "Overall Experience"
    series #series {
      value: count(surveyDataset_SA.response:OA1)
      label: "Overall Experience"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:OA1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    description: "Overall, I was able to find and understand the information I needed to pick an insurance plan."
  }
  label: "SA_OA1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #SA_OA3_stacked_bar {
  widget chart #SA_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "SALES - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_SA.response:OA3)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }
  label: "SA_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #SA_PA_stacked_bar {
  label: "SA_PA stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #SA_PA_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Provider Availability"
    series #series {
      value: count(ProviderAvailability:value)
      label: "Provider Availability"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: ProviderAvailability:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #SA_PA_Components_stacked_bar {
  label: "SA_PA Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #SA_PA_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Provider Availability Components"
    series #series {
      value: count(ProviderAvailability:value)
      label: "Provider Availability"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: ProviderAvailability:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: ProviderAvailability:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #SA_PA_grid {
  label: "SA_PA grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #SA_PA_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(ProviderAvailability:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_SA:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: ProviderAvailability:field
      showLabel: false
      totalLabel: "Provider Availability"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #SA_PA_trend_line {
  widget chart #SAtrendchart {
    cardCorners: '20px'
    label: "What are SALES - Provider Availability scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Provider Availability"
      value: average(numeric(ProviderAvailability:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Existing PCP in network"
      value: average(numeric(surveyDataset_SA:SA_PA2))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Existing spec in network"
      value: average(numeric(surveyDataset_SA:SA_PA4))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Hospital/facility in network"
      value: average(numeric(surveyDataset_SA:SA_PA5))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "PCP local"
      value: average(numeric(surveyDataset_SA:SA_PA6))
      format: OneDecimalNumberFormatter
    }
    series #series_6 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Spec local"
      value: average(numeric(surveyDataset_SA:SA_PA7))
      format: OneDecimalNumberFormatter
    }
    series #series_7 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Finding provider(s) that meet certain characteristics"
      value: average(numeric(surveyDataset_SA:SA_PA8))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "SALES - PA Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "SA_PA trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_PA_KDA_Correlation {
  label: "SA_PA KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #SA_OA2_PA_keyDriversWidget {
    cardCorners: '20px'
    label: "Provider Availability Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_SA:OA2
    independentVariables: surveyDataset_SA:SA_PA2, surveyDataset_SA:SA_PA4, surveyDataset_SA:SA_PA5, surveyDataset_SA:SA_PA6, surveyDataset_SA:SA_PA7, surveyDataset_SA:SA_PA8
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 62
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #SA_PA_Drilldown {
  label: "SA_PA Drilldown"
  widget canvas #SA_PA_SectionDrilldown_divider_canvasWidget {
    label: "SA_PA Section Drilldowns Divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "52px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Provider Availability Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #SA_PA_DrilldownResponses_canvasWidget {
    cardCorners: '20px'
    label: "SA_PA Drilldown responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "46px"
        left: "18px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "38px"
        left: "70px"
      }
      area #area_3 {
        position: "absolute"
        top: "169px"
        left: "70px"
      }
      area #area_4 {
        position: "absolute"
        top: "178px"
        left: "18px"
      }
      area #area_5 {
        position: "absolute"
        top: "288px"
        left: "70px"
      }
      area #area_6 {
        position: "absolute"
        top: "46px"
        left: "370px"
      }
      area #area_7 {
        position: "absolute"
        top: "38px"
        left: "422px"
      }
      area #area_8 {
        position: "absolute"
        top: "169px"
        left: "422px"
      }
      area #area_9 {
        position: "absolute"
        top: "178px"
        left: "370px"
      }
      area #area_10 {
        position: "absolute"
        top: "288px"
        left: "422px"
      }
      area #area_11 {
        position: "absolute"
        top: "80px"
        left: "720px"
      }
      area #area_12 {
        position: "absolute"
        top: "72px"
        left: "772px"
      }
      area #area_15 {
        position: "absolute"
        top: "288px"
        left: "772px"
      }
      area #area_16 {
        position: "absolute"
        top: "80px"
        left: "1097px"
      }
      area #area_17 {
        position: "absolute"
        top: "72px"
        left: "1149px"
      }
      area #area_20 {
        position: "absolute"
        top: "288px"
        left: "1123px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "70px"
      }
      area #area_19 {
        position: "absolute"
        top: "0px"
        left: "397px"
      }
      area #area_21 {
        position: "absolute"
        top: "0px"
        left: "741px"
      }
      area #area_22 {
        position: "absolute"
        top: "0px"
        left: "1094px"
      }
      background: #ffffff
    }
    tile value #valueTile {
      areaId: "area"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "Disagreed that it was easy to find out if their current PCP was covered and                                            "
      areaId: "area_2"
      style #style {
        width: "214px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile text #SA_PA2_B2BforDD_textTile {
      value: "Disagreed that it was easy to find a PCP nearby"
      areaId: "area_3"
      style #style {
        width: "248px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile value #valueTile_2 {
      areaId: "area_4"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_3 {
      value: "Among those who disagreed"
      areaId: "area_5"
      style #style {
        fontSize: 24
        width: "169px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PA_PCP_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PA4)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_4 {
      value: "Disagreed that it was easy to find out if their current specialist was covered and                                            "
      areaId: "area_7"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_5 {
      value: "Disagreed that it was easy to find a specialist nearby"
      areaId: "area_8"
      style #style {
        fontSize: 24
        width: "225px"
        height: "34px"
        color: #02253b
      }
    }
    tile value #valueTile_4 {
      areaId: "area_9"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PA7)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_6 {
      value: "Among those who disagreed"
      areaId: "area_10"
      style #style {
        fontSize: 24
        width: "167px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PA_Specialist_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PA5)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_7 {
      value: "Disagreed that it was easy to find out if their preferred hospital was covered                                            "
      areaId: "area_12"
      style #style {
        fontSize: 24
        width: "236px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_9 {
      value: "Among those who disagreed"
      areaId: "area_15"
      style #style {
        fontSize: 24
        width: "168px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PA_Hospital_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_7 {
      areaId: "area_16"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PA8)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_10 {
      value: "Disagreed that it was easy to find provider(s) that met personal preferences and needs                                         "
      areaId: "area_17"
      style #style {
        fontSize: 24
        width: "206px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_12 {
      value: "Among those who disagreed"
      areaId: "area_20"
      style #style {
        fontSize: 24
        width: "168px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PA_PersonalPreferrence_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #textTile_11 {
      value: "Finding a PCP"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_13 {
      value: "Finding a Specialist"
      areaId: "area_19"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_14 {
      value: "Finding a preferred Hospital"
      areaId: "area_21"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "231px"
        height: "47px"
      }
    }
    tile text #textTile_15 {
      value: "Finding preferred providers"
      areaId: "area_22"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "226px"
        height: "82px"
      }
    }
    cardTransparent: true
  }
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_PA_PCP_Drilldown {
  label: "SA_PA_PCP_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Where members tried to find information about a PCP"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_SA:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_SA:SA_DD1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Where members tried to find information about a PCP"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD1.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD1.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PA2_PA6_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about a PCP"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
        mode: "clustered"
      }
      value: count(surveyDataset_SA:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_SA:SA_DD2
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about a PCP"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD2.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD2.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "Members were able to eventually find out information about PCPs"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD3
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about PCPs"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD4)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD4
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
    description: "Select one."
  }
  widget comments #commentsWidget_3 {
    cardCorners: '20px'
    label: "Where members eventually found information about PCPs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD4.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD4.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_PA_Specialist_Drilldown {
  label: "SA_PA_Specialist_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Where members tried to find information about a Specialist"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_SA:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_SA:SA_DD5
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Where members tried to find information about a Specialist"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD5.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD5.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PA4_PA7_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about a Specialist"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
        mode: "clustered"
      }
      value: count(surveyDataset_SA:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_SA:SA_DD6
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_5 {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about a Specialist"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD6.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD6.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "Members were able to eventually find out information about Specialists"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD7
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about Specialists"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD8)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD8
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
    description: "Select one."
  }
  widget comments #commentsWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about Specialists"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD8.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD8.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_PA_Hospital_Drilldown {
  label: "SA_PA_Hospital_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Where members tried to find information about their preferred hospital"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_SA:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_SA:SA_DD9
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Where members tried to find information about their preferred hospital"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD9.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD9.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PA5_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about their preferred hospital"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD10
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_7 {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about their preferred hospital"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD10.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD10.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "Members were able to eventually find out information about their preferred hospital"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD11
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about preferred hospitals"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD12)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD12
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget_8 {
    cardCorners: '20px'
    label: "Where members eventually found information about preferred hospitals"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD12.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD12.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_PA_PersonalPreferrence_Drilldown {
  label: "SA_PA_PersonalPreferrence_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Where members tried to find information about preferred providers"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD13
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Where members tried to find information about their preferred providers"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD13.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD13.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PA8_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about preferred providers"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD14
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_9 {
    cardCorners: '20px'
    label: "Why members said it was difficult to find information about their preferred providers"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD14.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD14.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "Members were able to eventually find out information about preferred providers"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD15
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about preferred providers"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD16)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD16
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget_10 {
    cardCorners: '20px'
    label: "Where members eventually found information about preferred providers"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD16.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD16.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_RX_stacked_bar {
  label: "SA_RX stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #SA_RX_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rx Availability"
    series #series {
      value: count(RxAvailability:value)
      label: "Rx Availability"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: RxAvailability:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #SA_RX_Components_stacked_bar {
  label: "SA_RX Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #SA_RX_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rx Availability Components"
    series #series {
      value: count(RxAvailability:value)
      label: "Rx Availability"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 42
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: RxAvailability:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: RxAvailability:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #SA_RX_grid {
  label: "SA_RX grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #SA_PA_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(RxAvailability:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_SA:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: RxAvailability:field
      showLabel: false
      totalLabel: "Rx Availability"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #SA_RX_trend_line {
  widget chart #SAtrendchart {
    cardCorners: '20px'
    label: "What are SALES - Pharmacy/Rx Availability scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Pharmacy/Rx Availability"
      value: average(numeric(RxAvailability:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Preferred pharmacy local"
      value: average(numeric(surveyDataset_SA:SA_RX2))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Mail order Rx available"
      value: average(numeric(surveyDataset_SA:SA_RX3))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Other local pharmacy"
      value: average(numeric(surveyDataset_SA:SA_RX4))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rx cost"
      value: average(numeric(surveyDataset_SA:SA_RX5))
      format: OneDecimalNumberFormatter
    }
    description: "SALES - RX Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "SA_RX trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_RX_KDA_Correlation {
  label: "SA_RX KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #SA_OA2_RX_keyDriversWidget {
    cardCorners: '20px'
    label: "Rx Availability Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_SA:OA2
    independentVariables: surveyDataset_SA:SA_RX2, surveyDataset_SA:SA_RX6, surveyDataset_SA:SA_RX3, surveyDataset_SA:SA_RX4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    importanceLimit: 0
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #SA_RX_Drilldown {
  label: "SA_RX Drilldown"
  widget canvas #SA_RX_SectionDrilldown_divider_canvasWidget {
    label: "SALES Rx Section Drilldowns divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "52px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Rx Availability Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #SA_RX_DrilldownResponses_canvasWidget {
    label: "SA_RX Drilldown responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "72px"
        left: "46px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "63px"
        left: "98px"
      }
      area #area_3 {
        position: "absolute"
        top: "186px"
        left: "98px"
      }
      area #area_4 {
        position: "absolute"
        top: "195px"
        left: "46px"
      }
      area #area_5 {
        position: "absolute"
        top: "288px"
        left: "98px"
      }
      area #area_6 {
        position: "absolute"
        top: "72px"
        left: "572px"
      }
      area #area_7 {
        position: "absolute"
        top: "63px"
        left: "624px"
      }
      area #area_10 {
        position: "absolute"
        top: "288px"
        left: "624px"
      }
      area #area_11 {
        position: "absolute"
        top: "80px"
        left: "1031px"
      }
      area #area_12 {
        position: "absolute"
        top: "72px"
        left: "1083px"
      }
      area #area_15 {
        position: "absolute"
        top: "288px"
        left: "1083px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "58px"
      }
      area #area_19 {
        position: "absolute"
        top: "0px"
        left: "561px"
      }
      area #area_21 {
        position: "absolute"
        top: "0px"
        left: "1052px"
      }
    }
    tile value #valueTile {
      areaId: "area"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_RX2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        background: "#ffffff"
        borderRadius: "13.6px"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #SA_B2BforRXDD_textTile_1 {
      value: "Disagreed that it was easy to find out if their preferred pharmacy was covered and                                            "
      areaId: "area_2"
      style #style {
        width: "257px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile text #SA_B2BforRXDD_textTile_2 {
      value: "Disagreed that it was easy to find a pharmacy nearby"
      areaId: "area_3"
      style #style {
        width: "248px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile value #valueTile_2 {
      areaId: "area_4"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_RX4)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #SA_B2BforRXDD_textTile_3 {
      value: "Among those who disagreed"
      areaId: "area_5"
      style #style {
        fontSize: 24
        width: "169px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_RX_PreferredPharmacy_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_RX3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #SA_B2BforRXDD_textTile_4 {
      value: "Disagreed that it was easy to find out if they could get their prescription medicines by mail order                                 "
      areaId: "area_7"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #SA_B2BforRXDD_textTile_5 {
      value: "Among those who disagreed"
      areaId: "area_10"
      style #style {
        fontSize: 24
        width: "167px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_RX_MailOrder_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #SA_B2BforRXDD_textTile_6 {
      areaId: "area_11"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_RX5)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #SA_B2BforRXDD_textTile_7 {
      value: "Disagreed that they were able to understand what their current medications would cost                                            "
      areaId: "area_12"
      style #style {
        fontSize: 24
        width: "236px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #SA_B2BforRXDD_textTile_8 {
      value: "Among those who disagreed"
      areaId: "area_15"
      style #style {
        fontSize: 24
        width: "168px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_RX_MedicationCost_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #SA_B2BforRXDD_textTile_9 {
      value: "Finding a preferred pharmacy"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "250px"
        height: "79px"
      }
    }
    tile text #SA_B2BforRXDD_textTile_10 {
      value: "Finding mail-order information"
      areaId: "area_19"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "294px"
        height: "85px"
      }
    }
    tile text #SA_B2BforRXDD_textTile_11 {
      value: "Finding medication costs"
      areaId: "area_21"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "231px"
        height: "47px"
      }
    }
  }
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_RX_PreferredPharmacy_Drilldown {
  label: "SA_RX_PreferredPharmacy_Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about their preferred pharmacy"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD17
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    label: "Where members tried to find information about their preferred pharmacy"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD17.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD17.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_RX_PreferredPharmacy_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about a preferred pharmacy"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD18
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about their preferred pharmacy"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD18.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD18.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about their preferred pharmacy"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD3
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about preferred pharmacies"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD20)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD20
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget_3 {
    label: "Where members eventually found information about preferred pharmacies"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      comment: surveyDataset_SA:SA_DD20.98$other
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD20.98$other != ""
      }
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_RX_MailOrder_Drilldown {
  label: "SA_RX_MailOrder_Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about their mail order medications"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD21
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    label: "Where members tried to find information about their mail order medications"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD21.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD21.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_RX_MailOrder_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about mail order medications"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD22
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about their mail order medications"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD22.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD22.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about their mail order medications"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD23
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about mail order medications"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD24)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD24
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget_3 {
    label: "Where members eventually found information about mail order medications"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      comment: surveyDataset_SA:SA_DD24.98$other
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD24.98$other != ""
      }
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_RX_MedicationCost_Drilldown {
  label: "SA_RX_MedicationCost_Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about their current medication cost"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD25
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    label: "Where members tried to find information about their current medication cost"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD25.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD25.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_RX_RxCost_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about current medication cost"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD26
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about their current medication cost"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD26.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD26.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about their current medication cost"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD27
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about current medication cost"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD28)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD28
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget_3 {
    label: "Where members eventually found information about current medication cost"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      comment: surveyDataset_SA:SA_DD28.98$other
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD28.98$other != ""
      }
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_PC_stacked_bar {
  label: "SA_PC stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #SA_PC_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Premium/Coverages"
    series #series {
      value: count(PremiumCoverages:value)
      label: "Premium/Coverages"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: PremiumCoverages:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #SA_PC_Components_stacked_bar {
  label: "SA_PC Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #SA_PC_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Premium/Coverages Components"
    series #series {
      value: count(PremiumCoverages:value)
      label: "Premium/Coverages"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 42
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: PremiumCoverages:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: PremiumCoverages:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #SA_PC_grid {
  label: "SA_PC grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #SA_PA_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(PremiumCoverages:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_SA:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: PremiumCoverages:field
      showLabel: false
      totalLabel: "Premium/Coverages"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #SA_PC_trend_line {
  widget chart #SAtrendchart {
    cardCorners: '20px'
    label: "What are SALES - Premium/Coverages scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Premium/Coverages"
      value: average(numeric(PremiumCoverages:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Understand cost of plan"
      value: average(numeric(surveyDataset_SA:SA_PC1))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Understand cost of care"
      value: average(numeric(surveyDataset_SA:SA_PC2))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Covered services"
      value: average(numeric(surveyDataset_SA:SA_PC3))
      format: OneDecimalNumberFormatter
    }
    description: "SALES - PC Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "SA_PC trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_PC_SB_KDA_Correlation {
  label: "SA_PC_SB KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #SA_OA2_PC_keyDriversWidget {
    cardCorners: '20px'
    label: "Premium/Coverages and Supplemental Benefits Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_SA:OA2
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    independentVariables: surveyDataset_SA:SA_PC1, surveyDataset_SA:SA_PC2, surveyDataset_SA:SA_PC3, surveyDataset_SA:SA_SB1
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #SA_PC_Drilldown {
  label: "SA_PC Drilldown"
  widget canvas #SA_PC_SectionDrilldown_divider_canvasWidget {
    label: "SALES PC Section Drilldowns Divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "52px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Premium/Coverages Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #SA_PC_DrilldownResponses_canvasWidget {
    label: "SA_PC Drilldown Responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "97px"
        left: "18px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "89px"
        left: "70px"
      }
      area #area_5 {
        position: "absolute"
        top: "288px"
        left: "70px"
      }
      area #area_7 {
        position: "absolute"
        top: "97px"
        left: "586px"
      }
      area #area_10 {
        position: "absolute"
        top: "288px"
        left: "601px"
      }
      area #area_11 {
        position: "absolute"
        top: "105px"
        left: "534px"
      }
      area #area_16 {
        position: "absolute"
        top: "97px"
        left: "1071px"
      }
      area #area_17 {
        position: "absolute"
        top: "89px"
        left: "1123px"
      }
      area #area_20 {
        position: "absolute"
        top: "288px"
        left: "1123px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "70px"
      }
      area #area_19 {
        position: "absolute"
        top: "0px"
        left: "576px"
      }
      area #area_22 {
        position: "absolute"
        top: "0px"
        left: "1094px"
      }
    }
    tile value #valueTile {
      areaId: "area"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PC1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        background: "#ffffff"
        borderRadius: "13.6px"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "Disagreed that they were able to find monthly health insurance cost info                                            "
      areaId: "area_2"
      style #style {
        width: "214px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile text #textTile_3 {
      value: "Among those who disagreed"
      areaId: "area_5"
      style #style {
        fontSize: 24
        width: "169px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PC_PremiumCosts_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #textTile_4 {
      value: "Disagreed that they were able to understand what the costs for medical care would be                                            "
      areaId: "area_7"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_6 {
      value: "Among those who disagreed"
      areaId: "area_10"
      style #style {
        fontSize: 24
        width: "167px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PC_MedicalCareCost_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PC2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile value #valueTile_7 {
      areaId: "area_16"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_PC3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_10 {
      value: "Disagreed that they were able to find info about covered care and services                        "
      areaId: "area_17"
      style #style {
        fontSize: 24
        width: "206px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_12 {
      value: "Among those who disagreed"
      areaId: "area_20"
      style #style {
        fontSize: 24
        width: "168px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_PC_CareService_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #textTile_11 {
      value: "Finding premium cost"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_13 {
      value: "Finding OOP cost"
      areaId: "area_19"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_15 {
      value: "Finding care/service coverage info"
      areaId: "area_22"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "226px"
        height: "110px"
      }
    }
  }
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_PC_PremiumCosts_Drilldown {
  label: "SA_PC_PremiumCosts_Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about premium costs"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD29
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    label: "Where members tried to find information about their premium costs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD29.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD29.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PC1_PremCost_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about premium costs"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD30
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about their premium costs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD30.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD30.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about premium costs"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD31
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about premium costs"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD32)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD32
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget_3 {
    label: "Where members eventually found information about premium costs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD32.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD32.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_PC_MedicalCareCost_Drilldown {
  label: "SA_PC_MedicalCareCost_Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about medical care costs"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD33
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_3 {
    label: "Where members tried to find information about medical care costs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD33.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD33.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PC2_HCCost_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about medical care costs"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD34
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about medical care costs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD34.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD34.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about medical care costs"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD35
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about medical care costs"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD36)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD36
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget {
    label: "Where members eventually found information about medical care costs"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD36.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD36.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_PC_CareService_Drilldown {
  label: "SA_PC_CareService_Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about covered care and services"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD37
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_3 {
    label: "Where members tried to find information about covered care and services"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD37.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD37.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_PC3_CareSvc_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about covered care and services"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD38
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about covered care and services"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD38.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD38.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about covered care and services"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD39
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about covered care and services"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD40)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD40
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget {
    label: "Where members eventually found information about covered care and services"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD40.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD40.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_SB1_stacked_bar {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "Supplemental Benefits"
    series #series {
      value: count(surveyDataset_SA.response:SA_SB1)
      label: "Supplemental Benefits"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_SB1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
  }
  label: "SA_SB1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #SA_SB_grid {
  label: "SA_SB grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #SA_PA_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(surveyDataset_SA:SA_SB1))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_SA:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
    row #row {
      label: "Supplemental Benefits"
    }
  }
}





page #SA_SB_trend_line {
  widget chart #SAtrendchart {
    cardCorners: '20px'
    label: "What are SALES - Supplemental Benefits scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Supplemental Benefits"
      value: average(numeric(surveyDataset_SA:SA_SB1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_SA:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
    }
    description: "SALES - SB Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "SA_SB trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_SB_Drilldown_divider {
  label: "SA_SB Drilldown"
  widget canvas #SA_SB_SectionDrilldown_divider_canvasWidget {
    label: "SA_SB Section Drilldowns divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "52px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "SALES Supplemental Benefits Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #SA_SB_Drilldwown_canvasWidget {
    label: "SA_SB Drilldown"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "115px"
        left: "518px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "98px"
        left: "588px"
      }
      area #area_5 {
        position: "absolute"
        top: "288px"
        left: "600px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "506px"
      }
    }
    tile value #valueTile {
      areaId: "area"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_SA.response:SA_SB1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        background: "#ffffff"
        borderRadius: "13.6px"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "Disagreed that they were able to understand what additional benefits would be covered                                            "
      areaId: "area_2"
      style #style {
        width: "214px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile text #textTile_3 {
      value: "Among those who disagreed"
      areaId: "area_5"
      style #style {
        fontSize: 24
        width: "169px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "SA_SB_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #textTile_11 {
      value: "Finding covered additional benefits"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
  }
  hide: false
  modal: true
  modalSize: "large"
}





page #SA_SB_Drilldown {
  label: "SA_SB Drilldown charts"
  widget chart #chartWidget_5 {
    label: "Where members tried to find information about covered additional benefits"
    series #series {
      chart bar #barChart {
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD41
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_3 {
    label: "Where members tried to find information about covered additional benefits"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD41.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD41.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #SA_SB1_Drilldown_chartWidget {
    label: "Why members said it was difficult to find information about covered additional benefits"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
      }
      value: count(surveyDataset_SA:respid)
      percentOver: "categories"
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    category cutByMulti #cutCategory {
      value: surveyDataset_SA:SA_DD42
      valuePosition: outer
      sortOrder: descending
      sortBy: "series"
    }
    size: medium
    legend: "none"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    label: "Why members said it was difficult to find information about covered additional benefits"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD42.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD42.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  widget chart #chartWidget_4 {
    label: "Members were able to eventually find out information about covered additional benefits"
    series #series {
      value: surveyDataset_SA:numberOfResponses()
      format: PercentOneDecimalFormatter
      percentOver: "categories"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    chart pie #pieChart {
    }
    legend: "rightTop"
    category cut #cutCategory {
      value: surveyDataset_SA:SA_DD43
    }
  }
  widget chart #chartWidget_6 {
    cardCorners: '20px'
    label: "Where members eventually found information about covered additional benefits"
    series #series {
      value: count(surveyDataset_SA.response:SA_DD44)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_SA:SA_DD44
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    layout: "vertical"
  }
  widget comments #commentsWidget {
    label: "Where members eventually found information about covered additional benefits"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:SA_DD44.98$other != ""
      }
      comment: surveyDataset_SA:SA_DD44.98$other
    }
    size: "medium"
    table: surveyDataset_SA:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}





page #SA_Comments {
  label: "SA Comments"
  hide: false
  modal: true
  modalSize: "large"
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "What did members have to say about their SALES experience?"
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_SA:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_SA:OA2 != ""
      }
      comment: surveyDataset_SA:OA2
    }
    size: large
    table: surveyDataset_SA:
    cardBackground: #ffffff
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_SA.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #valueColumn {
      label: "Gender"
      value: surveyDataset_SA.response:ITGENDER
      align: center
      enableColumnFilter: true
    }
  }


}




















page #ENROLL {





  label: "ENROLLMENT"
}





page #ONBOARDING {





  label: "ONBOARDING"
}





page #FINDING_DRS {





  label: "FINDING CARE"
}










page #BENEFITS_USAGE {
  widget canvas #BENEFITS_USAGE_canvasWidget {
    label: "BENEFITS USAGE report links"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
      area #area_3 {
        position: "absolute"
        top: "6px"
        left: "555px"
      }
      area #area_5 {
        position: "absolute"
        top: "6px"
        left: "828px"
      }
      area #area_6 {
        position: "absolute"
        top: "6px"
        left: "1100px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Links to BENEFITS USAGE Components"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
    tile text #textTile_2 {
      value: "ACCESS TO CARE"
      areaId: "area_3"
      style #style {
        width: "259px"
        height: "31px"
        textAlign: "center"
        border: "solid medium #ffffff"
        borderRadius: "13.6px"
        padding: "1px 8px 8px 8px"
        fontWeight: "bold"
        background: "#ffffff"
        fontSize: 18
      }
      navigateTo: "ACCESS_TO_CARE"
      navigateOptions: "same_tab"
    }
  }
  label: "BENEFITS USAGE"
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1
}





page #ACCESS_TO_CARE {





  label: "BENEFITS USAGE - ACCESS TO CARE"
  widget canvas #AC_KPI_scores_divider {
    label: "AC type of care divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE : What type of care was this visit for? "
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #copy_of_AC_KPIScores_tabs_divider {
    label: "AC type of care tabs divider"
    container: container position {
      width: 1368px
      height: "55px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "338px"
      }
      area #area_5 {
        top: "17px"
        left: "139px"
        position: "absolute"
      }
      area #area_6 {
        top: "17px"
        left: "477px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "140px"
      }
      area #area_12 {
        position: "absolute"
        top: "35px"
        left: "478px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Urgent care"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #textTile_3 {
      value: "Routine care"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: PercentageOfAnswers(surveyDataset_AC.response:AC_MA1, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: PercentageOfAnswers(surveyDataset_AC.response:AC_MA1, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_AC.response:AC_MA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_AC.response:AC_MA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget canvas #copy_of_AC_KPI_scores_divider {
    label: "Copy of AC KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #AC_KPIScores_tabs_divider {
    label: "AC KPI scores tabs divider"
    container: container position {
      width: 1368px
      height: "55px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "845px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1183px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "7px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "6px"
        left: "1326px"
      }
      area #area_10 {
        top: "32px"
        left: "309px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "832px"
      }
      area #area_12 {
        position: "absolute"
        top: "34px"
        left: "1170px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Overall Experience"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #AC_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_AC.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: average(numeric(surveyDataset_AC:OA1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_AC:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "AC_OA2_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "AC_OA1_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "AC_OA3_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_AC.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_AC.response:OA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_AC.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #AC_NPS_trendchart {
    cardCorners: '20px'
    label: "How is ACCESS TO CARE NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_AC.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #AC_KPI_trendchart {
    cardCorners: '20px'
    label: "How are ACCESS TO CARE KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Overall Experience with ACCESS TO CARE"
      value: average(numeric(surveyDataset_AC:OA1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_AC:OA3))
      format: OneDecimalNumberFormatter
    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #AC_KeyDrivers_divider {
    label: "AC Key Drivers of KPIs divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE Key Drivers of KPIs"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget keyDrivers #AC_OA2_keyDriversWidget {
    cardCorners: '20px'
    label: "NPS"
    size: medium
    dependentVariable: surveyDataset_AC:OA2
    independentVariables: surveyDataset_AC:AC_MA2, surveyDataset_AC:AC_MA3, surveyDataset_AC:AC_MA4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.89
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #AC_OA1_keyDriversWidget {
    cardCorners: '20px'
    label: "Overall Experience"
    size: small
    dependentVariable: surveyDataset_AC:OA1
    independentVariables: surveyDataset_AC:AC_MA2, surveyDataset_AC:AC_MA3, surveyDataset_AC:AC_MA4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.89
    importanceLimit: 0.03
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #AC_OA3_keyDriversWidget {
    cardCorners: '20px'
    label: "Rating of Health Plan"
    size: small
    dependentVariable: surveyDataset_AC:OA3
    independentVariables: surveyDataset_AC:AC_MA2, surveyDataset_AC:AC_MA3, surveyDataset_AC:AC_MA4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.89
    importanceLimit: 0.03
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget canvas #AC_Section_scores_divider {
    label: "AC Section scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE Section scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #AC_SectionScores_tabs_divider {
    label: "AC Section scores tabs divider"
    container: container position {
      width: 1368px
      height: "59px"
      background: rgba(255, 255, 255, 0)
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "140px"
        position: "absolute"
      }
      area #area_9 {
        position: "absolute"
        top: "35px"
        left: "140px"
      }
      area #area_13 {
        position: "absolute"
        top: "6px"
        left: "297px"
      }
    }
    cardTransparent: true

    tile text #AC_MA_textTile {
      value: "Making Appointments"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Making Appointments"
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "Making Appointments"
      value: average(numeric(MakingAppts:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_9"
      label: "Making Appointments"
      value: count(surveyDataset_AC:respid, numeric(surveyDataset_AC:AC_MA2) >= 0 OR numeric(surveyDataset_AC:AC_MA3) >= 0 OR numeric(surveyDataset_AC:AC_MA4) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }

    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_13"
      style #style {
        width: "34px"
      }
      navigateTo: "AC_MA_stacked_bar"
      navigateOptions: "same_tab"
    }
  }
  widget chart #AC_SectionScore_trendchart {
    cardCorners: '20px'
    label: "How are ACCESS TO CARE Section scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Making Appointments"
      value: average(numeric(MakingAppts:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }
    }
    description: ""
    size: large
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #AC_ScoreComparison_divider {
    label: "AC Score Comparison divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_AC:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_AC:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_AC:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_AC:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_AC:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_AC:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_AC:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_AC.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_AC:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Making Appointments Composite'
        value: {
          qid: MakingAppts:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of contacting provider'
        value: {
          qid: surveyDataset_AC:AC_MA2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of scheduling appointment'
        value: {
          qid: surveyDataset_AC:AC_MA3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Received appointment as soon as needed'
        value: {
          qid: surveyDataset_AC:AC_MA4
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: false
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget chart #AC_ScoreComparison_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_AC:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_AC:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_AC:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_AC:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_AC:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_AC:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_AC:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
      item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_AC.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
      item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_AC:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Making Appointments Composite'
        value: {
          qid: MakingAppts:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of contacting provider'
        value: {
          qid: surveyDataset_AC:AC_MA2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Ease of scheduling appointment'
        value: {
          qid: surveyDataset_AC:AC_MA3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Received appointment as soon as needed'
        value: {
          qid: surveyDataset_AC:AC_MA4
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #AC_SectionCompoenentScores_divider {
    label: "AC Section and Component Scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE Section and Component Scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget headline #AC_MA_Dial {
    cardCorners: '20px'
    label: "Making Appointments"
    tile gauge #gaugeTile {
      value: average(numeric(MakingAppts:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "AC_MA_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"

    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_22__row {
        value: surveyDataset_AC:Dial__gridTile_22__variable$field

      }
      cell #Dial__gridTile_22__column__cell {
        value: average(numeric(surveyDataset_AC:Dial__gridTile_22__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_22__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_22__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_22__column {
        hide: false
      }
      sort rows #Dial__gridTile_22__sort {
        sortBy: "/Dial__gridTile_22__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_22__row
        column: @Dial__gridTile_22__column
        cell: @Dial__gridTile_22__column__cell
        sort: @Dial__gridTile_22__sort
        variable: @Dial__gridTile_22__variable
        chartColumn: @Dial__gridTile_22__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "AC_MA_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "AC_MA_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "AC_MA_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button.png"
      padding: true
      navigateTo: "AC_MA_Drilldown"
      navigateOptions: "same_tab"
    }
  }
  widget canvas #AC_Comment_divider {
    label: "AC Comment divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall ACCESS TO CARE experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please provide any additional comments."
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_AC:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_AC:OA4 != ""
      }
      comment: surveyDataset_AC:OA4
    }
    size: large
    table: surveyDataset_AC:
    cardBackground: #ffffff
    column value #AC_OA1_valueColumn {
      label: "Overall Experience Response"
      value: surveyDataset_AC.response:OA1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_AC.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #AC_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_AC.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #AC_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_AC.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #AC_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_AC.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #AC_Response_divider {
    label: "AC Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #AC_surveyMetricsWidget {
    cardCorners: '20px'
    label: "ACCESS TO CARE Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_AC
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1
  hide: true
  modal: false
}




page #AC_OA2_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "ACCESS TO CARE NPS"
    series #series {
      value: count(surveyDataset_AC.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_AC:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "On a scale of 0 to 10, how likely are you to recommend this health plan to a friend or a colleague?"
    layout: "vertical"
  }
  widget headline #AC_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_AC.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_AC.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #AC_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_AC.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_AC.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #AC_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_AC.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_AC.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "AC_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #AC_OA1_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "Overall Satisfaction with Access to Care"
    series #series {
      value: count(surveyDataset_AC.response:OA1)
      label: "Overall Experience"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_AC:OA1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    description: "Overall, I was satisfied with my ability to get appointments for the care I needed."
  }
  label: "AC_OA1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #AC_OA3_stacked_bar {
  widget chart #AC_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "ACCESS TO CARE - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_AC.response:OA3)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_AC:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }
  label: "AC_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}




page #AC_MA_stacked_bar {
  label: "AC_MA stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #AC_MA_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Making Appointments"
    series #series {
      value: count(MakingAppts:value)
      label: "Making Appointments"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: MakingAppts:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #AC_MA_Components_stacked_bar {
  label: "AC_MA Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #AC_MA_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Making Appointments Components"
    series #series {
      value: count(MakingAppts:value)
      label: "Making Appointments"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: MakingAppts:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: MakingAppts:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #AC_MA_grid {
  label: "AC_MA grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #AC_MA_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(MakingAppts:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_AC:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: MakingAppts:field
      showLabel: false
      totalLabel: "Making Appointments"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #AC_MA_trend_line {
  widget chart #ACtrendchart {
    cardCorners: '20px'
    label: "What are ACCESS TO CARE - Making Appointments scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false

      }
      label: "Making Appointments"
      value: average(numeric(MakingAppts:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_AC:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Ease of contacting provider"
      value: average(numeric(surveyDataset_AC:AC_MA2))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Ease of scheduling appointment"
      value: average(numeric(surveyDataset_AC:AC_MA3))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Seen in adequate time"
      value: average(numeric(surveyDataset_AC:AC_MA4))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "ACCESS TO CARE - MA Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "AC_MA trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #AC_MA_KDA_Correlation {
  label: "AC_MA KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #AC_OA2_MA_keyDriversWidget {
    cardCorners: '20px'
    label: "Making Appointments Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_AC:OA2
    independentVariables: surveyDataset_AC:AC_MA2, surveyDataset_AC:AC_MA3, surveyDataset_AC:AC_MA4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 49.89
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #AC_MA_Drilldown {
  label: "AC_MA Drilldown"
  widget canvas #AC_MA_SectionDrilldown_divider_canvasWidget {
    label: "AC_MA Section Drilldowns Divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "52px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "ACCESS TO CARE Making Appointments Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #AC_MA_Drilldown {
    label: "AC_MA Drilldown Responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "97px"
        left: "240px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "89px"
        left: "292px"
      }
      area #area_5 {
        position: "absolute"
        top: "288px"
        left: "292px"
      }
      area #area_16 {
        position: "absolute"
        top: "97px"
        left: "735px"
      }
      area #area_17 {
        position: "absolute"
        top: "89px"
        left: "787px"
      }
      area #area_20 {
        position: "absolute"
        top: "288px"
        left: "787px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "243px"
      }
      area #area_22 {
        position: "absolute"
        top: "0px"
        left: "758px"
      }
    }
    tile value #valueTile {
      areaId: "area"
      label: "Contacting provider"
      value: bottom2percent(surveyDataset_AC.response:AC_MA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        background: "#ffffff"
        borderRadius: "13.6px"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "Disagreed that it was easy to contact their provider"
      areaId: "area_2"
      style #style {
        width: "214px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile text #textTile_3 {
      value: "Among those who disagreed"
      areaId: "area_5"
      style #style {
        fontSize: 24
        width: "169px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "AC_MA_Contact_Drilldown"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_7 {
      areaId: "area_16"
      label: "Scheduling appointments"
      value: bottom2percent(surveyDataset_AC.response:AC_MA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_10 {
      value: "Disagreed that it was easy to schedule an appointment with their provider"
      areaId: "area_17"
      style #style {
        fontSize: 24
        width: "206px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_12 {
      value: "Among those who disagreed"
      areaId: "area_20"
      style #style {
        fontSize: 24
        width: "168px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "AC_MA_Appt_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #textTile_11 {
      value: "Contact provider"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_15 {
      value: "Scheduling appointments"
      areaId: "area_22"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "226px"
        height: "110px"
      }
    }
  }
  hide: false
  modal: true
  modalSize: "large"
}





page #AC_MA_Contact_Drilldown {
  label: "AC_MA_Contact_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "What were the difficulties that members experienced when trying to contact their provider?"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_AC:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_AC:AC_DD1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Other things members had difficulty with when trying to contact their provider"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_AC:AC_DD1.98$other != ""
      }
      comment: surveyDataset_AC:AC_DD1.98$other
    }
    size: "medium"
    table: surveyDataset_AC:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}




page #AC_MA_Appt_Drilldown {
  label: "AC_MA_Appt_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Difficulties experienced when trying to schedule an appointment with their provider?"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_AC:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_AC:AC_DD2
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Other difficulties with when trying to schedule an appointment with their provider"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_AC:AC_DD2.98$other != ""
      }
      comment: surveyDataset_AC:AC_DD2.98$other
    }
    size: "medium"
    table: surveyDataset_AC:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}










page #RX_MGMT {





  label: "RX MANAGEMENT"

  widget canvas #RXMGMT_REPORT_LINKS {
    label: "RX MGMT report links"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
      area #area_3 {
        position: "absolute"
        top: "6px"
        left: "555px"
      }
      area #area_5 {
        position: "absolute"
        top: "6px"
        left: "828px"
      }
      area #area_6 {
        position: "absolute"
        top: "6px"
        left: "1100px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Links to RX MANAGEMENT Components"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
    tile text #textTile_2 {
      value: "RX PREAUTHORIZATION"
      areaId: "area_3"
      style #style {
        width: "259px"
        height: "31px"
        textAlign: "center"
        border: "solid medium #ffffff"
        borderRadius: "13.6px"
        padding: "1px 8px 8px 8px"
        fontWeight: "bold"
        background: "#ffffff"
        fontSize: 18
      }
      navigateTo: "RX_MGMT_RXPREAUTH"
      navigateOptions: "same_tab"
    }
    tile text #textTile_3 {
      value: "GETTING PRESCRIPTIONS"
      areaId: "area_5"
      style #style {
        width: "259px"
        height: "31px"
        textAlign: "center"
        border: "solid medium #ffffff"
        borderRadius: "13.6px"
        padding: "1px 8px 8px 8px"
        fontWeight: "bold"
        background: "#ffffff"
        fontSize: 18
      }
      navigateTo: "RX_MGMT_GETTINGRX"
      navigateOptions: "same_tab"
    }
    tile text #textTile_4 {
      value: "RX CONCIERGE SERVICES"
      areaId: "area_6"
      style #style {
        width: "259px"
        height: "31px"
        textAlign: "center"
        border: "solid medium #ffffff"
        borderRadius: "13.6px"
        padding: "1px 8px 8px 8px"
        fontWeight: "bold"
        background: "#ffffff"
        fontSize: 18
      }
      navigateTo: "RX_MGMT_CONRX"
      navigateOptions: "same_tab"
    }
  }
  widget canvas #RXMGMT_KPI_scores_divider {
    label: "RX MGMT KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX MANAGEMENT KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #RXMGMT_KPIScores_tabs_divider {
    label: "RXMGMT KPI scores tabs divider"
    container: container position {
      width: 1368px
      height: "55px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "838px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1176px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "7px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "6px"
        left: "1326px"
      }
      area #area_10 {
        top: "32px"
        left: "309px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "832px"
      }
      area #area_12 {
        position: "absolute"
        top: "34px"
        left: "1170px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Overall Satisfaction"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #RXMGMT_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_RXCombo.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: average(numeric(surveyDataset_RXCombo:OA1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_RXCombo:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "RXMGMT_NPS_stacked"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "RXMGMT_OA1_stacked"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "RXMGMT_OA3_stacked"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_RXCombo.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_RXCombo.response:OA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_RXCombo.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #RP_NPS_trendchart {
    cardCorners: '20px'
    label: "How is RX MANAGEMENT NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_RXCombo.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_RXCombo:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_RXCombo:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #RXMGMT_KPI_trendchart {
    cardCorners: '20px'
    label: "How are RX MANAGEMENT KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Overall Experience with RX MANAGEMENT"
      value: average(numeric(surveyDataset_RXCombo:OA1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_RXCombo:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_RXCombo:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_RXCombo:OA3))
      format: OneDecimalNumberFormatter
    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }

  widget canvas #RXMGMT_ScoreComparison_divider {
    label: "RXMGMT Score Comparison divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX MANAGEMENT Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RXCombo:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RXCombo:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RXCombo:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RXCombo:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RXCombo:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RXCombo:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_RXCombo:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_RXCombo.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_RXCombo:OA3
          target: 48
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10
    }
  }
  widget chart #RXMGMT_ScoreComparison_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RXCombo:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RXCombo:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RXCombo:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RXCombo:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RXCombo:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RXCombo:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_RXCombo:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_RXCombo.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_RXCombo:OA3
          target: 48
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #RXMGMT_Comment_divider {
    label: "RXMGMT Comment divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall RX MANAGEMENT experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please provide any additional comments."
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_RXCombo:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_RXCombo:OA4 != ""
      }
      comment: surveyDataset_RXCombo:OA4
    }
    size: large
    table: surveyDataset_RXCombo:
    cardBackground: #ffffff
    column value #RP_OA1_valueColumn {
      label: "Overall Experience Response"
      value: surveyDataset_RXCombo.response:OA1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_RXCombo.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #RXMGMT_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_RXCombo.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #RXMGMT_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_RXCombo.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #RXMGMT_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_RXCombo.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #RXMGMT_Response_divider {
    label: "RXMGMT Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX MANAGEMENT Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #RXMGMT_surveyMetricsWidget {
    cardCorners: '20px'
    label: "RX MANAGEMENT Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_RXCombo
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4
}
page #RXMGMT_NPS_stacked {
  widget chart #RXMGMT_NPS_stacked_chartWidget {
    cardCorners: '20px'
    label: "RX MANAGEMENT NPS"
    series #series {
      value: count(surveyDataset_RXCombo.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_RXCombo:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "On a scale of 0 to 10, how likely are you to recommend this health plan to a friend or a colleague?"
    layout: "vertical"
  }
  widget headline #RXMGMT_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_RXCombo.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_RXCombo.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #RXMGMT_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_RXCombo.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_RXCombo.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #RXMGMT_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_RXCombo.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_RXCombo.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "RXMGMT_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}
page #RXMGMT_OA1_stacked {
  widget chart #RXMGMT_OA1_stacked_chartWidget {
    cardCorners: '20px'
    label: "Overall Satisfaction with Rx Management"
    series #series {
      value: count(surveyDataset_RXCombo.response:OA1)
      label: "Overall Experience"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_RXCombo:OA1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    description: "Overall Satisfaction"
  }
  label: "RXMGMT_OA1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}
page #RXMGMT_OA3_stacked {
  widget chart #RXMGMT_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "RX MANAGEMENT - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_RXCombo.response:OA3)
      label: "RHP"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_RXCombo:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }
  label: "RXMGMT_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #RX_MGMT_RXPREAUTH {





  label: "RX MANAGMENT - RX PREAUTHORIZATION"
  widget canvas #RP_PREAUTH_NOTE_scores_divider {
    label: "RP rcvd preauth note divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #RP_PREAUTH_NOTE_tabs_divider {
    label: "RP preauth note tabs divider"
    container: container position {
      width: 1368px
      height: "171px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "36px"
        left: "0px"
      }
      area #area_4 {
        position: "absolute"
        top: "36px"
        left: "338px"
      }
      area #area_5 {
        top: "44px"
        left: "139px"
        position: "absolute"
      }
      area #area_6 {
        top: "46px"
        left: "481px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "64px"
        left: "140px"
      }
      area #area_12 {
        position: "absolute"
        top: "65px"
        left: "478px"
      }
      area #area_7 {
        position: "absolute"
        top: "36px"
        left: "676px"
      }
      area #area_8 {
        position: "absolute"
        top: "36px"
        left: "1014px"
      }
      area #area_9 {
        position: "absolute"
        top: "46px"
        left: "815px"
      }
      area #area_10 {
        position: "absolute"
        top: "47px"
        left: "1158px"
      }
      area #area_13 {
        position: "absolute"
        top: "65px"
        left: "816px"
      }
      area #area_14 {
        position: "absolute"
        top: "65px"
        left: "1154px"
      }
      area #area_15 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_16 {
        position: "absolute"
        top: "0px"
        left: "676px"
      }
      area #area_17 {
        position: "absolute"
        top: "112px"
        left: "338px"
      }
      area #area_18 {
        position: "absolute"
        top: "113px"
        left: "676px"
      }
      area #area_19 {
        position: "absolute"
        top: "132px"
        left: "477px"
      }
      area #area_20 {
        position: "absolute"
        top: "132px"
        left: "819px"
      }
      area #area_21 {
        position: "absolute"
        top: "151px"
        left: "478px"
      }
      area #area_22 {
        position: "absolute"
        top: "149px"
        left: "816px"
      }
      area #area_23 {
        position: "absolute"
        top: "89px"
        left: "0px"
      }
      area #area_24 {
        position: "absolute"
        top: "145px"
        left: "564px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Yes"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile text #textTile_3 {
      value: "No"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "68px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "RP PA2 Yes"
      value: PercentageOfAnswers(surveyDataset_RP.response:RP_PA1, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
        width: "60px"
        height: "40px"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RP PA2 No"
      value: PercentageOfAnswers(surveyDataset_RP.response:RP_PA1, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "RP PA2 BASE"
      value: count(surveyDataset_RP.response:RP_PA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "RP PA2 BASE"
      value: count(surveyDataset_RP.response:RP_PA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_4 {
      value: "Yes"
      areaId: "area_7"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile text #textTile_5 {
      value: "No"
      areaId: "area_8"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile value #valueTile_7 {
      areaId: "area_9"
      label: "RP PA2 Yes"
      value: PercentageOfAnswers(surveyDataset_RP.response:RP_PA2, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_8 {
      areaId: "area_10"
      label: "RP PA2 No"
      value: PercentageOfAnswers(surveyDataset_RP.response:RP_PA2, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_9 {
      areaId: "area_13"
      label: "RP PA2 BASE"
      value: count(surveyDataset_RP.response:RP_PA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_10 {
      areaId: "area_14"
      label: "RP PA2 BASE"
      value: count(surveyDataset_RP.response:RP_PA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_6 {
      value: "Medications required preauthorization"
      areaId: "area_15"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "676px"
        height: "35px"
        textAlign: "center"
        border: "solid thin rgba(210, 255, 255, 0.14)"
        borderRadius: "0%"
        background: "#d2ffff"
      }
    }
    tile text #textTile_7 {
      value: "Received preauthorization notification"
      areaId: "area_16"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "676px"
        height: "35px"
        textAlign: "center"
        border: "solid thin rgba(210, 255, 255, 0.14)"
        borderRadius: "0%"
        background: "#d2ffff"
      }
    }
    tile text #textTile_8 {
      value: "Yes"
      areaId: "area_17"
      style #style {
        fontSize: 16
        width: "338px"
        height: "66px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "12px 8px 8px 8px"
      }
    }
    tile text #textTile_9 {
      value: "No"
      areaId: "area_18"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "65px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "12px 8px 8px 8px"
      }
    }
    tile value #valueTile_11 {
      areaId: "area_19"
      label: "RP PA2 Yes"
      value: PercentageOfAnswers(surveyDataset_RP.response:RP_PA4, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_12 {
      areaId: "area_20"
      label: "RP PA2 No"
      value: PercentageOfAnswers(surveyDataset_RP.response:RP_PA4, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_13 {
      areaId: "area_21"
      label: "RP PA2 BASE"
      value: count(surveyDataset_RP.response:RP_PA4)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_14 {
      areaId: "area_22"
      label: "RP PA2 BASE"
      value: count(surveyDataset_RP.response:RP_PA4)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_10 {
      value: "Medications preauthorization was denied"
      areaId: "area_23"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        color: #02253b
        width: "1352px"
        height: "35px"
        textAlign: "center"
        border: "solid thin rgba(210, 255, 255, 0.14)"
        borderRadius: "0%"
        background: "#d2ffff"
        fontWeight: "bold"
      }
    }
    tile text #textTile_11 {
      value: "(Use page filter to look deeper)"
      areaId: "area_24"
      style #style {
        fontSize: 12
        width: "224px"
        height: "25px"
        textAlign: "center"
        padding: "2px 8px 2px 8px"
      }
    }
  }
  widget canvas #RP_KPI_scores_divider {
    label: "RP KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #RP_KPIScores_tabs_divider {
    label: "RP KPI scores tabs divider"
    container: container position {
      width: 1368px
      height: "55px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "838px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1176px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "7px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "6px"
        left: "1326px"
      }
      area #area_10 {
        top: "32px"
        left: "309px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "832px"
      }
      area #area_12 {
        position: "absolute"
        top: "34px"
        left: "1170px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Overall Satisfaction"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #RP_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_RP.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: average(numeric(surveyDataset_RP:OA1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_RP:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "RP_OA2_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "RP_OA1_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "RP_OA3_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_RP.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_RP.response:OA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_RP.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #RP_NPS_trendchart {
    cardCorners: '20px'
    label: "How is RX PREAUTHORIZATION NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_RP.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #RP_KPI_trendchart {
    cardCorners: '20px'
    label: "How are RX PREAUTHORIZATION KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Overall Experience with RX PREAUTHORIZATION"
      value: average(numeric(surveyDataset_RP:OA1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_RP:OA3))
      format: OneDecimalNumberFormatter
    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #RP_KeyDrivers_divider {
    label: "RP Key Drivers of KPIs divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION Key Drivers of KPIs"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget keyDrivers #RP_OA2_keyDriversWidget {
    cardCorners: '20px'
    label: "NPS"
    size: medium
    dependentVariable: surveyDataset_RP:OA2
    independentVariables: surveyDataset_RP:RP_PA3, surveyDataset_RP:RP_PA6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: 0.02
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #RP_OA1_keyDriversWidget {
    cardCorners: '20px'
    label: "Overall Experience"
    size: small
    dependentVariable: surveyDataset_RP:OA1
    independentVariables: surveyDataset_RP:RP_PA3, surveyDataset_RP:RP_PA6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: -0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #RP_OA3_keyDriversWidget {
    cardCorners: '20px'
    label: "Rating of Health Plan"
    size: small
    dependentVariable: surveyDataset_RP:OA3
    independentVariables: surveyDataset_RP:RP_PA3, surveyDataset_RP:RP_PA6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget canvas #RP_Section_scores_divider {
    label: "RP Section scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION Section scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #RP_SectionScores_tabs_divider {
    label: "RP Section scores tabs divider"
    container: container position {
      width: 1368px
      height: "59px"
      background: rgba(255, 255, 255, 0)
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "140px"
        position: "absolute"
      }
      area #area_9 {
        position: "absolute"
        top: "35px"
        left: "140px"
      }
      area #area_13 {
        position: "absolute"
        top: "6px"
        left: "297px"
      }
    }
    cardTransparent: true

    tile text #RP_PA_textTile {
      value: "Rx Preauthorization"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Rx Preauthorization"
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "Rx Preauthorization"
      value: average(numeric(RXPreAuth:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_9"
      label: "Rx Preauthorization"
      value: count(surveyDataset_RP:respid, numeric(surveyDataset_RP:RP_PA3) >= 0 OR numeric(surveyDataset_RP:RP_PA6) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }

    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_13"
      style #style {
        width: "34px"
      }
      navigateTo: "RP_PA_stacked_bar"
      navigateOptions: "same_tab"
    }
  }
  widget chart #RP_SectionScore_trendchart {
    cardCorners: '20px'
    label: "How are RX PREAUTHORIZATION Section scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Rx Preauthorization"
      value: average(numeric(RXPreAuth:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }
    }
    description: ""
    size: large
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #RP_ScoreComparison_divider {
    label: "RP Score Comparison divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RP:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_RP:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_RP.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_RP:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx Preauthorization Composite'
        value: {
          qid: RXPreAuth:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of authorization'
        value: {
          qid: surveyDataset_RP:RP_PA3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Clarity of denial reason'
        value: {
          qid: surveyDataset_RP:RP_PA6
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10
    }
  }
  widget chart #RP_ScoreComparison_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RP:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_RP:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_RP.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_RP:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx Preauthorization Composite'
        value: {
          qid: RXPreAuth:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of authorization'
        value: {
          qid: surveyDataset_RP:RP_PA3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Clarity of denial reason'
        value: {
          qid: surveyDataset_RP:RP_PA6
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #RP_SectionCompoenentScores_divider {
    label: "RP Section and Component Scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION Section and Component Scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget headline #RP_PA_Dial {
    cardCorners: '20px'
    label: "Rx Preauthorization"
    tile gauge #gaugeTile {
      value: average(numeric(RXPreAuth:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "RP_PA_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"

    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_32__row {
        value: surveyDataset_RP:Dial__gridTile_32__variable$field

      }
      cell #Dial__gridTile_32__column__cell {
        value: average(numeric(surveyDataset_RP:Dial__gridTile_32__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_32__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_32__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_32__column {
        hide: false
      }
      sort rows #Dial__gridTile_32__sort {
        sortBy: "/Dial__gridTile_32__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_32__row
        column: @Dial__gridTile_32__column
        cell: @Dial__gridTile_32__column__cell
        sort: @Dial__gridTile_32__sort
        variable: @Dial__gridTile_32__variable
        chartColumn: @Dial__gridTile_32__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "RP_PA_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "RP_PA_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "RP_PA_KDA_Correlation"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button%20red.png"
      padding: true
      navigateTo: "RP_PA_Drilldown"
      navigateOptions: "same_tab"
    }
  }
  widget caseList #caseListWidget {
    label: "Case List"
    size: halfwidth
    navigateTo: ActionMgmt
  }
  widget caseList #copy_of_caseListWidget {
    label: "Copy of Case List"
    size: halfwidth
    navigateTo: ActionMgmt
  }
  widget canvas #RP_Comment_divider {
    label: "RP Comment divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall RX PREAUTHORIZATION experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please provide any additional comments."
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_RP:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_RP:OA4 != ""
      }
      comment: surveyDataset_RP:OA4
    }
    size: large
    table: surveyDataset_RP:
    cardBackground: #ffffff
    column value #RP_OA1_valueColumn {
      label: "Overall Experience Response"
      value: surveyDataset_RP.response:OA1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_RP.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #RP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_RP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #RP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_RP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #RP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_RP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #RP_Response_divider {
    label: "RP Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #RP_surveyMetricsWidget {
    cardCorners: '20px'
    label: "RX PREAUTHORIZATION Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_RP
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_CX_LOB, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_OA1
  hide: true
  modal: false
  widget caseDetailsSummary #caseDetailsSummaryWidget {
    label: "Case Details Summary"
    size: "large"
  }
}





page #RP_OA2_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "RX PREAUTHORIZATION NPS"
    series #series {
      value: count(surveyDataset_RP.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_RP:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "On a scale of 0 to 10, how likely are you to recommend this health plan to a friend or a colleague?"
    layout: "vertical"
  }
  widget headline #RP_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_RP.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_RP.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #RP_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_RP.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_RP.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #RP_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_RP.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_RP.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "RP_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #RP_OA1_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "Overall Satisfaction with Rx Preauthorization"
    series #series {
      value: count(surveyDataset_RP.response:OA1)
      label: "Overall Experience"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_RP:OA1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    description: "Overall, I was satisfied with my ability to get appointments for the care I needed."
  }
  label: "RP_OA1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #RP_OA3_stacked_bar {
  widget chart #RP_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "RX PREAUTHORIZATION - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_RP.response:OA3)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_RP:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }
  label: "RP_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}




page #RP_PA_stacked_bar {
  label: "RP_PA stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #RP_PA_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rx Preauthorization"
    series #series {
      value: count(RXPreAuth:value)
      label: "Rx Preauthorization"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: RXPreAuth:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #RP_PA_Components_stacked_bar {
  label: "RP_PA Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #RP_PA_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rx Preauthorization Components"
    series #series {
      value: count(RXPreAuth:value)
      label: "Rx Preauthorization"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: RXPreAuth:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: RXPreAuth:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #RP_PA_grid {
  label: "RP_PA grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #RP_PA_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(RXPreAuth:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_RP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: RXPreAuth:field
      showLabel: false
      totalLabel: "Rx Preauthorization"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #RP_PA_trend_line {
  widget chart #RPtrendchart {
    cardCorners: '20px'
    label: "What are RX PREAUTHORIZATION - Rx Preauthorization scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Rx Preauthorization"
      value: average(numeric(RXPreAuth:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_RP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Timeliness of authorization"
      value: average(numeric(surveyDataset_RP:RP_PA3))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Clarity of reason for denial"
      value: average(numeric(surveyDataset_RP:RP_PA6))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "RX PREAUTHORIZATION - PA Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "RP_PA trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #RP_PA_KDA_Correlation {
  label: "RP_PA KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #RP_OA2_PA_keyDriversWidget {
    cardCorners: '20px'
    label: "Rx Preauthorization Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_RP:OA2
    independentVariables: surveyDataset_RP:RP_PA3, surveyDataset_RP:RP_PA6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: 0.02
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}





page #RP_PA_Drilldown {
  label: "RP_PA Drilldown"
  widget canvas #RP_PA_SectionDrilldown_divider_canvasWidget {
    label: "RP_PA Section Drilldowns Divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "52px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX PREAUTHORIZATION Rx Preauthorizations Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #RP_PA_Drilldown {
    label: "RP_PA Drilldown Responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "97px"
        left: "240px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "89px"
        left: "292px"
      }
      area #area_5 {
        position: "absolute"
        top: "288px"
        left: "292px"
      }
      area #area_16 {
        position: "absolute"
        top: "97px"
        left: "548px"
      }
      area #area_17 {
        position: "absolute"
        top: "89px"
        left: "608px"
      }
      area #area_20 {
        position: "absolute"
        top: "288px"
        left: "600px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "524px"
      }
      area #area_22 {
        position: "absolute"
        top: "0px"
        left: "758px"
      }
    }
    tile value #valueTile_7 {
      areaId: "area_16"
      label: "Clarity of reason for denial"
      value: bottom2percent(surveyDataset_RP.response:RP_PA6)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_10 {
      value: "Disagreed that they understood the reason for denial"
      areaId: "area_17"
      style #style {
        fontSize: 24
        width: "206px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_12 {
      value: "Among those who disagreed"
      areaId: "area_20"
      style #style {
        fontSize: 24
        width: "168px"
        height: "89px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "RP_PA_Timeliness_Drilldown"
      navigateOptions: "same_tab"
    }
    tile text #textTile_11 {
      value: "Clarity of reason for denial"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
  }
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "How many members disagreed compared across categories? (Highest 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RP:ITMEMST
      }
    }
    series #series {
      chart bar #barChart {
        showBase: false
      }
      value: bottom2percent(surveyDataset_RP.response:RP_PA6)
      valuePosition: outer
      label: ""
      format: PercentOneDecimalFormatter
      colorFormat: Single_Red_Color_Bar
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 by percentage are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10
    }
    palette: Single_Red_Color_Bar
  }
  widget chart #chartWidget_2 {
    cardCorners: '20px'
    label: "How many members disagreed compared across categories? (Lowest 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RP:ITMEMST
      }
    }
    series #series {
      chart bar #barChart {
        showBase: false
      }
      value: bottom2percent(surveyDataset_RP.response:RP_PA6)
      valuePosition: outer
      label: ""
      format: PercentOneDecimalFormatter
      colorFormat: Single_Red_Color_Bar
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 by percentage are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
    palette: Single_Red_Color_Bar
  }
  hide: false
  modal: true
  modalSize: "large"
}





page #RP_PA_Timeliness_Drilldown {
  label: "RP_PA_Clarity_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Difficulties experienced when trying to undertand the medication denial reasons"
    series #series {
      chart bar #barChart {
        mode: "clustered"
        showBase: true
        showValue: true
      }
      value: count(surveyDataset_RP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_RP:RP_DD1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."

    cardShadow: true
  }
  widget chart #chartWidget_2 {
    cardCorners: '20px'
    label: "Difficulties experienced by category"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RP:ITMEMST
      }
    }
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_RP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_RP:RP_DD1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "horizontal"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: large
    legend: "bottomLeft"
    description: "Multiple responses allowed."
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10
    }
  }
  widget dataGrid #dataGridWidget_3 {
    label: "Difficulties experienced by category (sortable table)"
    size: "medium"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_RP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_RP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_RP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_RP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_RP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_RP:ITMEMST
      }
    }
    column cut #column {
      value: @selectorBackgroundVar1.selected
      label: "Percent selected"
      cell rowPercentage #cell {
        value: count(surveyDataset_RP:respid)
        view: comparativeStatisticView
      }
    }
    row cutByMulti #row {
      value: surveyDataset_RP:RP_DD1
      total: "none"
    }
    description: "Click next to category columns to sort."
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      target: count(surveyDataset_RP.response:RP_DD1)
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: gridDefaultValueColorFormatter
      backgroundColorFormatter: gridDefaultBackgroundColorFormatter
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Other things members had difficulty understanding the reasons for denial"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_RP:RP_DD1.98$other != ""
      }
      comment: surveyDataset_RP:RP_DD1.98$other
    }
    size: "medium"
    table: surveyDataset_RP:
    description: "Other ( please specify)"
  }
  hide: false
  modal: true
}




page #RX_MGMT_GETTINGRX {





  label: "RX MANAGEMENT - GETTING PRESCRIPTIONS"
  widget canvas #GP_KPI_scores_divider {
    label: "GP KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #GP_KPIScores_tabs_divider {
    label: "GP KPI scores tabs divider"
    container: container position {
      width: 1368px
      height: "53px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "838px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1176px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "7px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "6px"
        left: "1326px"
      }
      area #area_10 {
        top: "32px"
        left: "309px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "832px"
      }
      area #area_12 {
        position: "absolute"
        top: "34px"
        left: "1170px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Overall Rating of Drug Plan"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #GP_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_GP.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: average(numeric(surveyDataset_GP:OA1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_GP:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "GettingRx_NPS_stacked"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "GP_OA1_stacked"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "GP_OA3_stacked"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_GP.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_GP.response:OA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_GP.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #GP_NPS_trendchart {
    cardCorners: '20px'
    label: "How is GETTING PRESCRIPTIONS NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_GP.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #GP_KPI_trendchart {
    cardCorners: '20px'
    label: "How are GETTING PRESCRIPTIONS KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Overall Rating of Drug Plan"
      value: average(numeric(surveyDataset_GP:OA1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_GP:OA3))
      format: OneDecimalNumberFormatter
    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #GP_RETAIL_scores_divider {
    label: "GP got Rx from retail divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #canvasWidget_12 {
    label: "RP preauth note tabs divider"
    container: container position {
      width: 1368px
      height: "88px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "36px"
        left: "0px"
      }
      area #area_4 {
        position: "absolute"
        top: "36px"
        left: "338px"
      }
      area #area_5 {
        top: "44px"
        left: "139px"
        position: "absolute"
      }
      area #area_6 {
        top: "46px"
        left: "481px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "64px"
        left: "140px"
      }
      area #area_12 {
        position: "absolute"
        top: "65px"
        left: "478px"
      }
      area #area_7 {
        position: "absolute"
        top: "36px"
        left: "676px"
      }
      area #area_8 {
        position: "absolute"
        top: "36px"
        left: "1014px"
      }
      area #area_9 {
        position: "absolute"
        top: "46px"
        left: "815px"
      }
      area #area_10 {
        position: "absolute"
        top: "47px"
        left: "1158px"
      }
      area #area_13 {
        position: "absolute"
        top: "65px"
        left: "816px"
      }
      area #area_14 {
        position: "absolute"
        top: "65px"
        left: "1154px"
      }
      area #area_15 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_16 {
        position: "absolute"
        top: "0px"
        left: "676px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Yes"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile text #textTile_3 {
      value: "No"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "68px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "RP PA2 Yes"
      value: PercentageOfAnswers(surveyDataset_GP.response:GP_RX1, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
        width: "60px"
        height: "40px"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RP PA2 No"
      value: PercentageOfAnswers(surveyDataset_GP.response:GP_RX1, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "RP PA2 BASE"
      value: count(surveyDataset_GP.response:GP_RX1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "RP PA2 BASE"
      value: count(surveyDataset_GP.response:GP_RX1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_4 {
      value: "Yes"
      areaId: "area_7"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile text #textTile_5 {
      value: "No"
      areaId: "area_8"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile value #valueTile_7 {
      areaId: "area_9"
      label: "RP PA2 Yes"
      value: PercentageOfAnswers(surveyDataset_GP.response:GP_MX1, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_8 {
      areaId: "area_10"
      label: "RP PA2 No"
      value: PercentageOfAnswers(surveyDataset_GP.response:GP_MX1, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_9 {
      areaId: "area_13"
      label: "RP PA2 BASE"
      value: count(surveyDataset_GP.response:GP_MX1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_10 {
      areaId: "area_14"
      label: "RP PA2 BASE"
      value: count(surveyDataset_GP.response:GP_MX1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile text #textTile_6 {
      value: "Got Rx from local pharmacy"
      areaId: "area_15"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "676px"
        height: "35px"
        textAlign: "center"
        border: "solid thin rgba(210, 255, 255, 0.14)"
        borderRadius: "0%"
        background: "#d2ffff"
      }
    }
    tile text #textTile_7 {
      value: "Got Rx from mail order pharmacy"
      areaId: "area_16"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "676px"
        height: "35px"
        textAlign: "center"
        border: "solid thin rgba(210, 255, 255, 0.14)"
        borderRadius: "0%"
        background: "#d2ffff"
      }
    }
  }
  widget canvas #GP_KeyDrivers_divider {
    label: "GP Key Drivers of KPIs divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS Key Drivers of KPIs"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget keyDrivers #GP_OA2_keyDriversWidget {
    cardCorners: '20px'
    label: "NPS"
    size: medium
    dependentVariable: surveyDataset_GP:OA2
    independentVariables: surveyDataset_GP:GP_RX2, surveyDataset_GP:GP_RX3, surveyDataset_GP:GP_RX4, surveyDataset_GP:GP_RX5, surveyDataset_GP:GP_RX6, surveyDataset_GP:GP_MX2, surveyDataset_GP:GP_MX3, surveyDataset_GP:GP_MX4, surveyDataset_GP:GP_MX5, surveyDataset_GP:GP_MX6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 52.1
    importanceLimit: 0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #GP_OA1_keyDriversWidget {
    cardCorners: '20px'
    label: "Overall Experience"
    size: small
    dependentVariable: surveyDataset_GP:OA1
    independentVariables: surveyDataset_GP:GP_RX2, surveyDataset_GP:GP_RX3, surveyDataset_GP:GP_RX4, surveyDataset_GP:GP_RX5, surveyDataset_GP:GP_RX6, surveyDataset_GP:GP_MX2, surveyDataset_GP:GP_MX3, surveyDataset_GP:GP_MX4, surveyDataset_GP:GP_MX5, surveyDataset_GP:GP_MX6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 52.1
    importanceLimit: .01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #GP_OA3_keyDriversWidget {
    cardCorners: '20px'
    label: "Rating of Health Plan"
    size: small
    dependentVariable: surveyDataset_GP:OA3
    independentVariables: surveyDataset_GP:GP_RX2, surveyDataset_GP:GP_RX3, surveyDataset_GP:GP_RX4, surveyDataset_GP:GP_RX5, surveyDataset_GP:GP_RX6, surveyDataset_GP:GP_MX2, surveyDataset_GP:GP_MX3, surveyDataset_GP:GP_MX4, surveyDataset_GP:GP_MX5, surveyDataset_GP:GP_MX6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 52.1
    importanceLimit: 0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget canvas #GP_Section_scores_divider {
    label: "GP Section scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS Section scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #GP_SectionScores_tabs_divider {
    label: "GP Section scores tabs divider"
    container: container position {
      width: 1368px
      height: "59px"
      background: rgba(255, 255, 255, 0)
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "140px"
        position: "absolute"
      }
      area #area_9 {
        position: "absolute"
        top: "35px"
        left: "140px"
      }
      area #area_13 {
        position: "absolute"
        top: "6px"
        left: "297px"
      }
      area #area_5 {
        position: "absolute"
        top: "0px"
        left: "338px"
      }
      area #area_6 {
        position: "absolute"
        top: "22px"
        left: "478px"
      }
      area #area_7 {
        position: "absolute"
        top: "33px"
        left: "478px"
      }
      area #area_8 {
        position: "absolute"
        top: "6px"
        left: "635px"
      }
    }
    cardTransparent: true

    tile text #GP_RX_textTile {
      value: "Retail Rx"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Retail Rx"
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "Retail Order Rx"
      value: average(numeric(RetailRX:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_9"
      label: "Retail Rx"
      value: count(surveyDataset_GP:respid, numeric(surveyDataset_GP:GP_RX2) >= 0 OR numeric(surveyDataset_GP:GP_RX3) >= 0 OR numeric(surveyDataset_GP:GP_RX4) >= 0 OR numeric(surveyDataset_GP:GP_RX5) >= 0 OR numeric(surveyDataset_GP:GP_RX6) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }

    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_13"
      style #style {
        width: "34px"
      }
      navigateTo: "GP_RX_stacked"
      navigateOptions: "same_tab"
    }
    tile text #textTile_2 {
      value: "Mail Order Rx"
      areaId: "area_5"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Retail Rx"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "Retail Order Rx"
      value: average(numeric(MailRX:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_4 {
      areaId: "area_7"
      label: "Mail Rx"
      value: count(surveyDataset_GP:respid, numeric(surveyDataset_GP:GP_MX2) >= 0 OR numeric(surveyDataset_GP:GP_MX3) >= 0 OR numeric(surveyDataset_GP:GP_MX4) >= 0 OR numeric(surveyDataset_GP:GP_MX5) >= 0 OR numeric(surveyDataset_GP:GP_MX6) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "GP_RX_stacked_bar"
      navigateOptions: "same_tab"
    }
  }
  widget chart #GP_SectionScore_trendchart {
    cardCorners: '20px'
    label: "How are GETTING PRESCRIPTIONS Section scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Retail Rx "
      value: average(numeric(RetailRX:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Mail Order Rx"
      value: average(numeric(MailRX:value)) * 1.33
      format: OneDecimalNumberFormatter
    }
    description: ""
    size: large
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #GP_ScoreComparison_divider {
    label: "GP Score Comparison divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RETAIL RX Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_GP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_GP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_GP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_GP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_GP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_GP:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Rating of Drug Plan'
        value: {
          qid: surveyDataset_GP:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_GP.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_GP:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Retail Rx Composite'
        value: {
          qid: RetailRX:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of getting retail prescription'
        value: {
          qid: surveyDataset_GP:GP_RX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Local pharmacy was courteous and respectful'
        value: {
          qid: surveyDataset_GP:GP_RX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Local pharmacy was helpful/answered questions'
        value: {
          qid: surveyDataset_GP:GP_RX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Easy to get refills at local pharmacy'
        value: {
          qid: surveyDataset_GP:GP_RX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Satisfied with local pharmacy'
        value: {
          qid: surveyDataset_GP:GP_RX6
          target: 87
          removeEmptyRows: true          
        }
      },
      item {
        label: 'Mail Order Rx Composite'
        value: {
          qid: MailRX:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of getting mail order prescription'
        value: {
          qid: surveyDataset_GP:GP_MX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order pharmacy was courteous and respectful'
        value: {
          qid: surveyDataset_GP:GP_MX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order pharmacy was helpful/answered questions'
        value: {
          qid: surveyDataset_GP:GP_MX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Easy to get mail order refills'
        value: {
          qid: surveyDataset_GP:GP_MX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Satisfied with mail order pharmacy'
        value: {
          qid: surveyDataset_GP:GP_MX6
          target: 87
          removeEmptyRows: true 
        }                  
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10
    }
  }
  widget chart #GP_ScoreComparison_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_GP:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_GP:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_GP:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_GP:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_GP:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_GP:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Rating of Drug Plan'
        value: {
          qid: surveyDataset_GP:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_GP.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_GP:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Retail Rx Composite'
        value: {
          qid: RetailRX:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of getting retail prescription'
        value: {
          qid: surveyDataset_GP:GP_RX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Local pharmacy was courteous and respectful'
        value: {
          qid: surveyDataset_GP:GP_RX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Local pharmacy was helpful/answered questions'
        value: {
          qid: surveyDataset_GP:GP_RX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Easy to get refills at local pharmacy'
        value: {
          qid: surveyDataset_GP:GP_RX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Satisfied with local pharmacy'
        value: {
          qid: surveyDataset_GP:GP_RX6
          target: 87
          removeEmptyRows: true          
        }
      },
      item {
        label: 'Mail Order Rx Composite'
        value: {
          qid: MailRX:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Timeliness of getting mail order prescription'
        value: {
          qid: surveyDataset_GP:GP_MX2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order pharmacy was courteous and respectful'
        value: {
          qid: surveyDataset_GP:GP_MX3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Mail order pharmacy was helpful/answered questions'
        value: {
          qid: surveyDataset_GP:GP_MX4
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Easy to get mail order refills'
        value: {
          qid: surveyDataset_GP:GP_MX5
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Satisfied with mail order pharmacy'
        value: {
          qid: surveyDataset_GP:GP_MX6
          target: 87
          removeEmptyRows: true 
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #GP_SectionCompoenentScores_divider {
    label: "GP Section and Component Scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS Section and Component Scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget headline #GP_RX_Dial {
    cardCorners: '20px'
    label: "Retail Rx"
    tile gauge #gaugeTile {
      value: average(numeric(RetailRX:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "GP_RX_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"

    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_33__row {
        value: surveyDataset_GP:Dial__gridTile_33__variable$field

      }
      cell #Dial__gridTile_33__column__cell {
        value: average(numeric(surveyDataset_GP:Dial__gridTile_33__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_33__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_33__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_33__column {
        hide: false
      }
      sort rows #Dial__gridTile_33__sort {
        sortBy: "/Dial__gridTile_33__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_33__row
        column: @Dial__gridTile_33__column
        cell: @Dial__gridTile_33__column__cell
        sort: @Dial__gridTile_33__sort
        variable: @Dial__gridTile_33__variable
        chartColumn: @Dial__gridTile_33__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "GP_RX_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "GP_RX_trend"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "GP_RX_KDA"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button%20red.png"
      padding: true
      navigateTo: "page_131"
      navigateOptions: "same_tab"
    }
  }
  widget headline #GP_MX_Dial {
    cardCorners: '20px'
    label: "Mail Order Rx"
    tile gauge #gaugeTile {
      value: average(numeric(MailRX:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "GP_MX_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"

    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_34__row {
        value: surveyDataset_GP:Dial__gridTile_34__variable$field

      }
      cell #Dial__gridTile_34__column__cell {
        value: average(numeric(surveyDataset_GP:Dial__gridTile_34__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_34__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_34__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_34__column {
        hide: false
      }
      sort rows #Dial__gridTile_34__sort {
        sortBy: "/Dial__gridTile_34__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_34__row
        column: @Dial__gridTile_34__column
        cell: @Dial__gridTile_34__column__cell
        sort: @Dial__gridTile_34__sort
        variable: @Dial__gridTile_34__variable
        chartColumn: @Dial__gridTile_34__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "GP_MX_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "GP_MX_trend"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "GP_MX_KDA"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_4 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Drilldown%20button%20red.png"
      padding: true
      navigateTo: "page_132"
      navigateOptions: "same_tab"
    }
  }
  widget canvas #GP_Comment_divider {
    label: "GP Comment divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall GETTING PRESCRIPTIONS experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please provide any additional comments."
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_GP:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:OA4 != ""
      }
      comment: surveyDataset_GP:OA4
    }
    size: large
    table: surveyDataset_GP:
    cardBackground: #ffffff
    column value #RP_OA1_valueColumn {
      label: "Overall Experience Response"
      value: surveyDataset_GP.response:OA1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_GP.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #GP_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_GP.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #GP_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_GP.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #GP_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_GP.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #GP_Response_divider {
    label: "GP Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #GP_surveyMetricsWidget {
    cardCorners: '20px'
    label: "GETTING PRESCRIPTIONS Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_GP
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4, fromQuestionFilter_CX_OA1, fromQuestionFilter_CX_MEMST, fromQuestionFilter_CX_RACE, fromQuestionFilter_CX_GENDER, fromQuestionFilter_CX_CONTRACT, fromQuestionFilter_CX_PLAN, fromQuestionFilter_CX_LOB
  hide: true
  modal: false
}
page #GettingRx_NPS_stacked {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "GETTING PRESCRIPTIONS NPS"
    series #series {
      value: count(surveyDataset_GP.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_GP:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "On a scale of 0 to 10, how likely are you to recommend this health plan to a friend or a colleague?"
    layout: "vertical"
  }
  widget headline #GP_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_GP.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_GP.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #GP_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_GP.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_GP.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #GP_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_GP.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_GP.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "GP_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}
page #GP_OA1_stacked {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "Overall Rating of Drug Plan"
    series #series {
      value: count(surveyDataset_GP.response:OA1)
      label: "Overall Experience"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_GP:OA1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    description: "Overall, I am satisfied with my prescription drug benefits."
  }
  label: "GP_OA1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}
page #GP_OA3_stacked {
  widget chart #GP_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "GETTING PRESCRIPTIONS - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_GP.response:OA3)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_GP:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }
  label: "GP_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}
page #GP_RX_stacked {
  label: "GP_RX stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #GP_RX_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Retail Rx"
    series #series {
      value: count(RetailRX:value)
      label: "Retail Rx"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: RetailRX:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}
page #GP_RX_Components_stacked_bar {
  label: "GP_RX Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #GP_RX_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Retail Rx Components"
    series #series {
      value: count(RetailRX:value)
      label: "Retail Rx"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: RetailRX:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: RetailRX:field
    }
    chartMargin {
      left: 30
      right: 35
      top: 0
    }
  }
}
page #GP_RX_grid {
  label: "GP_RX grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #GP_RX_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(RetailRX:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_GP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: RetailRX:field
      showLabel: false
      totalLabel: "Retail Rx"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}
page #GP_RX_trend {
  widget chart #GPtrendchart {
    cardCorners: '20px'
    label: "What are GETTING PRESCRIPTIONS - Retail Rx scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Retail Rx"
      value: average(numeric(RetailRX:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Timeliness of getting retail prescription"
      value: average(numeric(surveyDataset_GP:GP_RX2))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Local pharmacy was courteous and respectful"
      value: average(numeric(surveyDataset_GP:GP_RX3))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Local pharmacy was helpful/answered questions"
      value: average(numeric(surveyDataset_GP:GP_RX4))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Easy to get refills at local pharmacy"
      value: average(numeric(surveyDataset_GP:GP_RX5))
      format: OneDecimalNumberFormatter
    }
    series #series_6 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Satisfied with local pharmacy"
      value: average(numeric(surveyDataset_GP:GP_RX6))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "GETTING PRESCRIPTIONS - RX Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "GP_RX trend line"
  hide: false
  modal: true
  modalSize: "large"
}
page #GP_RX_KDA {
  label: "GP_RX KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #GP_OA2_RX_keyDriversWidget {
    cardCorners: '20px'
    label: "Retail Pharmacy Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_GP:OA2
    independentVariables: surveyDataset_GP:GP_RX2, surveyDataset_GP:GP_RX3, surveyDataset_GP:GP_RX4, surveyDataset_GP:GP_RX5, surveyDataset_GP:GP_RX6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 52.09
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}
page #page_131 {
  label: "GP_RX Drilldown"
  widget canvas #GP_RX_SectionDrilldown_divider_canvasWidget {
    label: "GP_RX Section Drilldowns Divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "61px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS Retail Rx Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #GP_RX_DrilldownResponses_canvasWidget {
    cardCorners: '20px'
    label: "GP_RX Drilldown responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "94px"
        left: "48px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "86px"
        left: "106px"
      }
      area #area_6 {
        position: "absolute"
        top: "86px"
        left: "328px"
      }
      area #area_7 {
        position: "absolute"
        top: "78px"
        left: "425px"
      }
      area #area_10 {
        position: "absolute"
        top: "294px"
        left: "329px"
      }
      area #area_11 {
        position: "absolute"
        top: "86px"
        left: "996px"
      }
      area #area_12 {
        position: "absolute"
        top: "78px"
        left: "1057px"
      }
      area #area_18 {
        position: "absolute"
        top: "8px"
        left: "116px"
      }
      area #area_19 {
        position: "absolute"
        top: "0px"
        left: "449px"
      }
      area #area_21 {
        position: "absolute"
        top: "0px"
        left: "1060px"
      }
      background: #ffffff
      area #area_13 {
        position: "absolute"
        top: "86px"
        left: "676px"
      }
      area #area_14 {
        position: "absolute"
        top: "79px"
        left: "745px"
      }
      area #area_17 {
        position: "absolute"
        top: "0px"
        left: "745px"
      }
    }
    tile value #valueTile {
      areaId: "area"
      label: "Got Rx as soon as needed"
      value: bottom2percent(surveyDataset_GP.response:GP_RX2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "Disagreed they got their meds from their local pharmacy as soon as needed                                            "
      areaId: "area_2"
      style #style {
        width: "214px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_GP.response:GP_RX3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_4 {
      value: "Disagreed that their local pharmacy treated them with courtesy and respect                                          "
      areaId: "area_7"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_6 {
      value: "Among those who disagreed"
      areaId: "area_10"
      style #style {
        fontSize: 24
        width: "746px"
        height: "44px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "GP_RX_Drilldown_charts"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_GP.response:GP_RX5)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_7 {
      value: "Disagreed that it was easy to get refills at their local pharmacy                                          "
      areaId: "area_12"
      style #style {
        fontSize: 24
        width: "236px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_11 {
      value: "Got Rx as soon
 as needed"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_13 {
      value: "Courtesy and
respect"
      areaId: "area_19"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_14 {
      value: "Getting Rx refills"
      areaId: "area_21"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "198px"
        height: "47px"
      }
    }
    cardTransparent: true
    tile value #valueTile_4 {
      areaId: "area_13"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_GP.response:GP_RX4)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_10 {
      value: "Disagreed that their local pharmacy was helpful in answering questions                                         "
      areaId: "area_14"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_15 {
      value: "Helpful answering questions"
      areaId: "area_17"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "228px"
        height: "110px"
      }
    }
  }
  hide: false
  modal: true
  modalSize: "large"
}
page #GP_RX_Drilldown_charts {
  label: "GP_RX_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Why getting Rx took longer than preferred"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_GP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_GP:GP_DD1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_4 {
    cardCorners: '20px'
    label: "Other reasons for not getting meds as soon as needed"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD1.98$other != ""
      }
      comment: surveyDataset_GP:GP_DD1.98$other
    }
    size: "medium"
    table: surveyDataset_GP:
    description: "Other (please specify)"
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "In what way was your local pharmacy not courteous of respectful?"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD2 != ""
      }
      comment: surveyDataset_GP:GP_DD2
    }
    size: "medium"
    table: surveyDataset_GP:
  }
  widget chart #SA_PA2_PA6_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Difficulties getting questions answered"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
        mode: "clustered"
      }
      value: count(surveyDataset_GP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_GP:GP_DD3
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    cardCorners: '20px'
    label: "Other difficulties with getting questions answered"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD3.98$other != ""
      }
      comment: surveyDataset_GP:GP_DD3.98$other
    }
    size: "medium"
    table: surveyDataset_GP:
    description: "Other (please specify)"
  }
  widget chart #GP_RX_RX5_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Difficulties getting refills"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
        mode: "clustered"
      }
      value: count(surveyDataset_GP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_GP:GP_DD4
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_3 {
    cardCorners: '20px'
    label: "Other difficulties with getting refills"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD4.98$other != ""
      }
      comment: surveyDataset_GP:GP_DD4.98$other
    }
    size: "medium"
    table: surveyDataset_GP:
  }
  hide: false
  modal: true
}

page #GP_MX_stacked_bar {
  label: "GP_MX stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #GP_MX_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Mail Order Rx"
    series #series {
      value: count(MailRX:value)
      label: "Mail Order Pharmacy"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: MailRX:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}
page #GP_MX_Components_stacked_bar {
  label: "GP_MX Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #GP_MX_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Mail Order Rx Components"
    series #series {
      value: count(MailRX:value)
      label: "Mail Order Pharmacy"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: MailRX:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: MailRX:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}
page #GP_MX_grid {
  label: "GP_MX grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #GP_MX_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(MailRX:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_GP:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: MailRX:field
      showLabel: false
      totalLabel: "Mail Order Pharmacy"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}
page #GP_MX_trend {
  widget chart #GPtrendchart {
    cardCorners: '20px'
    label: "What are GETTING PRESCRIPTIONS - Mail Order Pharmacy scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Mail Order Pharmacy"
      value: average(numeric(MailRX:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_GP:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Timeliness of getting mail order Rx"
      value: average(numeric(surveyDataset_GP:GP_MX2))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Mail order pharmacy was courteous and respectful"
      value: average(numeric(surveyDataset_GP:GP_MX3))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Mail order pharmacy was helpful/answered questions"
      value: average(numeric(surveyDataset_GP:GP_MX4))
      format: OneDecimalNumberFormatter
    }
    series #series_5 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Easy to get refills at mail order pharmacy"
      value: average(numeric(surveyDataset_GP:GP_MX5))
      format: OneDecimalNumberFormatter
    }
    series #series_6 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Satisfied with mail order pharmacy"
      value: average(numeric(surveyDataset_GP:GP_MX6))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "GETTING PRESCRIPTIONS - MX Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "GP_MX trend line"
  hide: false
  modal: true
  modalSize: "large"
}
page #GP_MX_KDA {
  label: "GP_MX KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #GP_OA2_MX_keyDriversWidget {
    cardCorners: '20px'
    label: "Mail Order Pharmacy Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_GP:OA2
    independentVariables: surveyDataset_GP:GP_MX2, surveyDataset_GP:GP_MX3, surveyDataset_GP:GP_MX4, surveyDataset_GP:GP_MX5, surveyDataset_GP:GP_MX6
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 52.09
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}
page #page_132 {
  label: "GP_MX Drilldown"
  widget canvas #GP_MX_SectionDrilldown_divider_canvasWidget {
    label: "GP_MX Section Drilldowns Divider"
    container: container position {
      width: 1368px
      height: "51px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "61px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "GETTING PRESCRIPTIONS Mail Order Rx Section Drilldown"
      areaId: "area_4"
      style #style {
        fontSize: 24
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #GP_MX_DrilldownResponses_canvasWidget {
    cardCorners: '20px'
    label: "GP_MX Drilldown responses"
    container: container position {
      width: 1368px
      height: "390px"
      area #area {
        top: "94px"
        left: "48px"
        position: "absolute"
      }
      area #area_2 {
        position: "absolute"
        top: "86px"
        left: "106px"
      }
      area #area_6 {
        position: "absolute"
        top: "86px"
        left: "328px"
      }
      area #area_7 {
        position: "absolute"
        top: "78px"
        left: "425px"
      }
      area #area_10 {
        position: "absolute"
        top: "294px"
        left: "329px"
      }
      area #area_11 {
        position: "absolute"
        top: "86px"
        left: "996px"
      }
      area #area_12 {
        position: "absolute"
        top: "78px"
        left: "1057px"
      }
      area #area_18 {
        position: "absolute"
        top: "8px"
        left: "116px"
      }
      area #area_19 {
        position: "absolute"
        top: "0px"
        left: "449px"
      }
      area #area_21 {
        position: "absolute"
        top: "0px"
        left: "1060px"
      }
      background: #ffffff
      area #area_13 {
        position: "absolute"
        top: "86px"
        left: "676px"
      }
      area #area_14 {
        position: "absolute"
        top: "77px"
        left: "745px"
      }
      area #area_17 {
        position: "absolute"
        top: "0px"
        left: "745px"
      }
    }
    tile value #valueTile {
      areaId: "area"
      label: "Got Rx as soon as needed"
      value: bottom2percent(surveyDataset_GP.response:GP_MX2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "Disagreed they got their mail order meds as soon as needed                                            "
      areaId: "area_2"
      style #style {
        width: "214px"
        height: "34px"
        color: #02253b
        fontSize: 24
      }
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "Courtesy and rspect"
      value: bottom2percent(surveyDataset_GP.response:GP_MX3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_4 {
      value: "Disagreed that the mail order pharmacy treated them with courtesy and respect                                          "
      areaId: "area_7"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_6 {
      value: "Among those who disagreed"
      areaId: "area_10"
      style #style {
        fontSize: 24
        width: "746px"
        height: "44px"
        textAlign: "center"
        padding: "8px 8px 8px 8px"
        background: "#D02541"
        borderRadius: "13.6px"
        color: #ffffff
      }
      label: "Among those who disagreed"
      navigateTo: "GP_MX_Drilldown_charts"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "Existing PCP in network"
      value: bottom2percent(surveyDataset_GP.response:GP_RX5)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_7 {
      value: "Disagreed that it was easy to get mail order refills                                          "
      areaId: "area_12"
      style #style {
        fontSize: 24
        width: "236px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_11 {
      value: "Got Rx as soon
 as needed"
      areaId: "area_18"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_13 {
      value: "Courtesy and
respect"
      areaId: "area_19"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
      }
    }
    tile text #textTile_14 {
      value: "Getting Rx refills"
      areaId: "area_21"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "198px"
        height: "47px"
      }
    }
    cardTransparent: true
    tile value #valueTile_4 {
      areaId: "area_13"
      label: "Helpful"
      value: bottom2percent(surveyDataset_GP.response:GP_MX4)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 24
        width: "52px"
        height: "34px"
        fontWeight: "bold"
        color: #02253b
      }
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile_10 {
      value: "Disagreed that the mail order pharmacy was helpful in answering questions                                         "
      areaId: "area_14"
      style #style {
        fontSize: 24
        width: "251px"
        height: "34px"
        color: #02253b
      }
    }
    tile text #textTile_15 {
      value: "Helpful answering questions"
      areaId: "area_17"
      style #style {
        fontSize: 24
        fontWeight: "bold"
        fontFamily: "Arial"
        textAlign: "center"
        textDecoration: "underline"
        color: #02253b
        width: "228px"
        height: "110px"
      }
    }
  }
  hide: false
  modal: true
  modalSize: "large"
}
page #GP_MX_Drilldown_charts {
  label: "GP_MX_Drilldown charts"
  widget chart #chartWidget_5 {
    cardCorners: '20px'
    label: "Why getting mail order Rx took longer than preferred"
    series #series {
      chart bar #barChart {
        mode: "clustered"
      }
      value: count(surveyDataset_GP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_GP:GP_DD5
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_4 {
    cardCorners: '20px'
    label: "Other reasons for not getting meds as soon as needed"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD5.98$other != ""
      }
      comment: surveyDataset_GP:GP_DD5.98$other
    }
    size: "medium"
    table: surveyDataset_GP:
    description: "Other (please specify)"
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "In what way was the mail order pharmacy not courteous or respectful?"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD6 != ""
      }
      comment: surveyDataset_GP:GP_DD6
    }
    size: "medium"
    table: surveyDataset_GP:
  }
  widget chart #SA_PA2_PA6_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Difficulties getting questions answered by mail order pharmacy"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
        mode: "clustered"
      }
      value: count(surveyDataset_GP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_GP:GP_DD7
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_2 {
    cardCorners: '20px'
    label: "Other difficulties with getting questions answered"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD7.98$other != ""
      }
      comment: surveyDataset_GP:GP_DD7.98$other
    }
    size: "medium"
    table: surveyDataset_GP:
    description: "Other (please specify)"
  }
  widget chart #GP_RX_RX5_Drilldown_chartWidget {
    cardCorners: '20px'
    label: "Difficulties getting mail order refills"
    series #series {
      chart bar #barChart {
        showBase: false
        showValue: true
        mode: "clustered"
      }
      value: count(surveyDataset_GP:respid)
      format: PercentOneDecimalFormatter
      palette: defaultColorPalette
      breakdownBy cutByMulti #cutBreakdownby {
        value: surveyDataset_GP:GP_DD8
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
      textSize: 100
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    layout: "vertical"
    removeEmptyCategories: true
    removeEmptySeries: false
    significanceTesting: false
    confidenceLevels: "95"
    size: medium
    legend: "rightTop"
    description: "Multiple responses allowed."
  }
  widget comments #commentsWidget_3 {
    cardCorners: '20px'
    label: "Other difficulties with getting refills"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Unlabeled Comment"
      filter expression #excludeBlankResponses {
        value: surveyDataset_GP:GP_DD8.98$other != ""
      }
      comment: surveyDataset_GP:GP_DD8.98$other
    }
    size: "medium"
    table: surveyDataset_GP:
  }
  hide: false
  modal: true
}

page #RX_MGMT_CONRX {





  label: "RX MANAGEMENT - RX CONCIERGE"
  widget canvas #CX_CONTACT_NOTE_scores_divider {
    label: "CX Contact note divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE - Contacted by the pharmacy team at your health insurance"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #CX_CONRX_NOTE_tabs_divider {
    label: "CX conrx note tabs divider"
    container: container position {
      width: 1368px
      height: "52px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "338px"
      }
      area #area_5 {
        top: "6px"
        left: "139px"
        position: "absolute"
      }
      area #area_6 {
        top: "8px"
        left: "477px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "26px"
        left: "140px"
      }
      area #area_12 {
        position: "absolute"
        top: "26px"
        left: "478px"
      }
      area #area_7 {
        position: "absolute"
        top: "0px"
        left: "676px"
      }
      area #area_8 {
        position: "absolute"
        top: "36px"
        left: "1014px"
      }
      area #area_9 {
        position: "absolute"
        top: "46px"
        left: "815px"
      }
      area #area_10 {
        position: "absolute"
        top: "47px"
        left: "1158px"
      }
      area #area_13 {
        position: "absolute"
        top: "65px"
        left: "816px"
      }
      area #area_14 {
        position: "absolute"
        top: "65px"
        left: "1154px"
      }
      area #area_15 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_16 {
        position: "absolute"
        top: "0px"
        left: "676px"
      }
      area #area_17 {
        position: "absolute"
        top: "0px"
        left: "338px"
      }
      area #area_18 {
        position: "absolute"
        top: "0px"
        left: "676px"
      }
      area #area_19 {
        position: "absolute"
        top: "132px"
        left: "477px"
      }
      area #area_20 {
        position: "absolute"
        top: "132px"
        left: "819px"
      }
      area #area_21 {
        position: "absolute"
        top: "151px"
        left: "478px"
      }
      area #area_22 {
        position: "absolute"
        top: "149px"
        left: "816px"
      }
      area #area_23 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_24 {
        position: "absolute"
        top: "145px"
        left: "564px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Yes"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile text #textTile_3 {
      value: "No"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "68px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
        padding: "3px 8px 8px 8px"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "CX CS1 Yes"
      value: PercentageOfAnswers(surveyDataset_CX.response:CX_CS1, "1")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
        width: "60px"
        height: "40px"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "CX CS1 No"
      value: PercentageOfAnswers(surveyDataset_CX.response:CX_CS1, "2")
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: PercentOneDecimalFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
        color: #000000
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "CX CS1 BASE"
      value: count(surveyDataset_CX.response:CX_CS1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "CX CS1 BASE"
      value: count(surveyDataset_CX.response:CX_CS1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget canvas #CX_KPI_scores_divider {
    label: "CX KPI scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE KPI scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #CX_KPIScores_tabs_divider {
    label: "CX KPI scores tabs divider"
    container: container position {
      width: 1368px
      height: "55px"
      background: rgba(255, 255, 255, 0)
      area #area {
        position: "absolute"
        top: "0px"
        left: "692px"
      }
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "309px"
        position: "absolute"
      }
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "1030px"
      }
      area #area_5 {
        top: "18px"
        left: "838px"
        position: "absolute"
      }
      area #area_6 {
        top: "18px"
        left: "1176px"
        position: "absolute"
      }
      area #area_7 {
        position: "absolute"
        top: "7px"
        left: "634px"
      }
      area #area_8 {
        position: "absolute"
        top: "7px"
        left: "988px"
      }
      area #area_9 {
        position: "absolute"
        top: "6px"
        left: "1326px"
      }
      area #area_10 {
        top: "32px"
        left: "309px"
        position: "absolute"
      }
      area #area_11 {
        position: "absolute"
        top: "34px"
        left: "832px"
      }
      area #area_12 {
        position: "absolute"
        top: "34px"
        left: "1170px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "Overall Satisfaction"
      areaId: "area"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile text #CX_NPS_textTile {
      value: "NPS"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "676px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "NPS"
      value: nps(surveyDataset_CX.response:OA2) * 100
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile text #textTile_3 {
      value: "Rating of Health Plan"
      areaId: "area_4"
      style #style {
        fontSize: 16
        fontFamily: "Trebuchet MS"
        fontWeight: "bold"
        color: #02253b
        width: "338px"
        height: "67px"
        textAlign: "center"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
    }
    tile value #valueTile_2 {
      areaId: "area_5"
      label: "Overall Experience"
      value: average(numeric(surveyDataset_CX:OA1))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile value #valueTile_3 {
      areaId: "area_6"
      label: "RHP"
      value: average(numeric(surveyDataset_CX:OA3))
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 16
        fontWeight: "bold"
      }
      view: valueDefaultView
      formatString: "{value}"
    }
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_7"
      style #style {
        width: "34px"
      }
      navigateTo: "CX_OA2_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_8"
      style #style {
        width: "34px"
      }
      navigateTo: "CX_OA1_Stacked_chartWidget"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_9"
      style #style {
        width: "34px"
      }
      navigateTo: "CX_OA3_stacked_bar"
      navigateOptions: "same_tab"
    }
    tile value #valueTile_4 {
      areaId: "area_10"
      label: "NPS"
      value: count(surveyDataset_CX.response:OA2)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_11"
      label: "NPS"
      value: count(surveyDataset_CX.response:OA1)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
    tile value #valueTile_6 {
      areaId: "area_12"
      label: "NPS"
      value: count(surveyDataset_CX.response:OA3)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }
  }
  widget chart #CX_NPS_trendchart {
    cardCorners: '20px'
    label: "How is RX CONCIERGE NPS trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "NPS"
      value: nps(surveyDataset_CX.response:OA2) * 100
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: -100
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget chart #CX_KPI_trendchart {
    cardCorners: '20px'
    label: "How are RX CONCIERGE KPI scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Overall Experience with RX CONCIERGE"
      value: average(numeric(surveyDataset_CX:OA1))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }

    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Rating of Health Plan"
      value: average(numeric(surveyDataset_CX:OA3))
      format: OneDecimalNumberFormatter
    }



    description: ""
    size: medium
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #CX_KeyDrivers_divider {
    label: "CX Key Drivers of KPIs divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE Key Drivers of KPIs"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget keyDrivers #CX_OA2_keyDriversWidget {
    cardCorners: '20px'
    label: "NPS"
    size: medium
    dependentVariable: surveyDataset_CX:OA2
    independentVariables: surveyDataset_CX:CX_CS2, surveyDataset_CX:CX_CS3, surveyDataset_CX:CX_CS4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: 0.02
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #CX_OA1_keyDriversWidget {
    cardCorners: '20px'
    label: "Overall Experience"
    size: small
    dependentVariable: surveyDataset_CX:OA1
    independentVariables: surveyDataset_CX:CX_CS2, surveyDataset_CX:CX_CS3, surveyDataset_CX:CX_CS4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: -0.01
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget keyDrivers #CX_OA3_keyDriversWidget {
    cardCorners: '20px'
    label: "Rating of Health Plan"
    size: small
    dependentVariable: surveyDataset_CX:OA3
    independentVariables: surveyDataset_CX:CX_CS2, surveyDataset_CX:CX_CS3, surveyDataset_CX:CX_CS4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: 0
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
    showModelDetails: true
    rSquaredLimit: 0.5
    defaultView: chart
  }
  widget canvas #CX_Section_scores_divider {
    label: "CX Section scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE Section scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget canvas #CX_SectionScores_tabs_divider {
    label: "CX Section scores tabs divider"
    container: container position {
      width: 1368px
      height: "59px"
      background: rgba(255, 255, 255, 0)
      area #area_2 {
        position: "absolute"
        top: "0px"
        left: "0px"
      }
      area #area_3 {
        top: "22px"
        left: "140px"
        position: "absolute"
      }
      area #area_9 {
        position: "absolute"
        top: "35px"
        left: "140px"
      }
      area #area_13 {
        position: "absolute"
        top: "6px"
        left: "297px"
      }
    }
    cardTransparent: true

    tile text #CX_CS_textTile {
      value: "Rx Concierge"
      areaId: "area_2"
      style #style {
        fontSize: 16
        width: "338px"
        height: "67px"
        textAlign: "center"
        fontFamily: "Trebuchet MS"
        color: #02253b
        fontWeight: "bold"
        border: "solid thin rgba(0, 0, 0, 0.14)"
        borderRadius: "13.6px"
        background: "#ffffff"
      }
      label: "Rx Concierge"
    }
    tile value #valueTile {
      areaId: "area_3"
      label: "Rx Concierge"
      value: average(numeric(ConRX:value))
      style #style {
        justifyContent: "center"
        alignItems: "center"
        width: "58px"
        height: "23px"
        fontSize: 16
        fontWeight: "bold"
      }
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      valueFormatter: OneDecimalNumberFormatter
    }
    tile value #valueTile_5 {
      areaId: "area_9"
      label: "Rx Concierge"
      value: count(surveyDataset_CX:respid, numeric(surveyDataset_CX:CX_CS2) >= 0 OR numeric(surveyDataset_CX:CX_CS3) >= 0 OR numeric(surveyDataset_CX:CX_CS4) >= 0)
      style #style {
        justifyContent: "center"
        alignItems: "center"
        fontSize: 11
        width: "58px"
        height: "30px"
      }
      valueFormatter: n_EqualsWithComma_baseFormatter
    }

    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/info%20dot.PNG"
      areaId: "area_13"
      style #style {
        width: "34px"
      }
      navigateTo: "CX_CS_stacked_bar"
      navigateOptions: "same_tab"
    }
  }
  widget chart #CX_SectionScore_trendchart {
    cardCorners: '20px'
    label: "How are RX CONCIERGE Section scores trending?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBaseInTooltip: true

      }
      label: "Rx Concierge"
      value: average(numeric(ConRX:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarMonth
            format: calendarMonthDefaultFormatter
          }
        }
      }
    }
    description: ""
    size: large
    legend: "bottomLeft"
    cardTransparent: false
    cardShadow: true
  }
  widget canvas #CX_ScoreComparison_divider {
    label: "CX Score Comparison divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE Score Comparison"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget chart #chartWidget_4 {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Top 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_CX:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_CX:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_CX:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_CX:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_CX:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_CX:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_CX:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_CX.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_CX:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx Concierge Composite'
        value: {
          qid: ConRX:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Helped save money'
        value: {
          qid: surveyDataset_CX:CX_CS2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Made sure taking meds correctly'
        value: {
          qid: surveyDataset_CX:CX_CS3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Helped coordinate with provider'
        value: {
          qid: surveyDataset_CX:CX_CS4
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Highest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: descending
      sortBy: "series"
      takeTop: 10
    }
  }
  widget chart #CX_ScoreComparison_chartWidget {
    cardCorners: '20px'
    label: "How do scores compare across categories? (Bottom 10)"
    select #selectorBackgroundVar1 {
      label: "Select a Category"
      options: item {
        label: 'Line of Business'
        value: surveyDataset_CX:ITLOB        
      },
      item {
        label: 'Plan Type'
        value: surveyDataset_CX:ITPLAN_TY
      },
      item {
        label: 'Contract'
        value: surveyDataset_CX:ITH_CONTRACT
      },
      item {
        label: 'Gender'
        value: surveyDataset_CX:ITGENDER
      },
      item {
        label: 'Race'
        value: surveyDataset_CX:ITRACE
      },
      item {
        label: 'Member State'
        value: surveyDataset_CX:ITMEMST
      }
    }
    select #selectorQuestion1 {
      label: "Select a Survey Measure"
      options: item {
        label: 'Overall Experience'
        value: {
          qid: surveyDataset_CX:OA1
          
          target: 77
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Likelihood to Recommend'
        value: {
          qid: surveyDataset_CX.response:OA2
          target: 48
          removeEmptyRows: true
        }
      },
       item { 
        label: 'Rating of Health Plan'
        value: {
          qid: surveyDataset_CX:OA3
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Rx Concierge Composite'
        value: {
          qid: ConRX:value
          target: 48
          removeEmptyRows: true
        }
      },
      item {
        label: 'Helped save money'
        value: {
          qid: surveyDataset_CX:CX_CS2
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Made sure taking meds correctly'
        value: {
          qid: surveyDataset_CX:CX_CS3
          target: 87
          removeEmptyRows: true
        }
      },
      item {
        label: 'Helped coordinate with provider'
        value: {
          qid: surveyDataset_CX:CX_CS4
          target: 87
          removeEmptyRows: true
        }
      }
    }
    series #series {
      chart bar #barChart {
        showBase: true
      }
      value: average(numeric(@selectorQuestion1.selected.qid))
      valuePosition: outer
      label: ""
      format: OneDecimalNumberFormatter
      colorFormat: SurveyResponseColorScaledMeanScoreFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    description: "For large categories -  Lowest 10 performers by score are shown."
    size: medium
    cardAlign: top
    removeEmptyCategories: true
    removeEmptySeries: true
    significanceTesting: true
    confidenceLevels: "95"
    legend: "none"
    category cut #cutCategory {
      value: @selectorBackgroundVar1.selected
      sortOrder: ascending
      sortBy: "series"
      takeTop: 10

    }
  }
  widget canvas #CX_SectionCompoenentScores_divider {
    label: "CX Section and Component Scores divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE Section and Component Scores"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget headline #CX_CS_Dial {
    cardCorners: '20px'
    label: "Rx Concierge"
    tile gauge #gaugeTile {
      value: average(numeric(ConRX:value))
      label: "Section Score"
      gaugeColorFormat: SurveyResponseColorScaledMeanScoreFormatter
      format: OneDecimalNumberFormatter
      min: 0
      showRange: true
      navigateTo: "CX_CS_Components_stacked_bar"
      navigateOptions: "same_tab"
      Composites trend #line {
      }
      target: 77
      max: 100
      aboveTargetLabel: "Above PG Benchmark"
      targetFormat: OneDecimalNumberFormatter
      belowTargetLabel: "Gap to PG Benchmark"
      atTargetLabel: "Meeting PG Benchmark"

    }
    cardTransparent: false
    cardShadow: false
    cardBackground: #ffffff
    cardText: #000000
    tile grid #gridTile {
      row cut #Dial__gridTile_35__row {
        value: surveyDataset_CX:Dial__gridTile_35__variable$field

      }
      cell #Dial__gridTile_35__column__cell {
        value: average(numeric(surveyDataset_CX:Dial__gridTile_35__variable$value))
        format: OneDecimalNumberFormatter
      }
      column #Dial__gridTile_35__chartColumn {
        width: "auto"
        cell microchart #microchartCell {
          value: @Dial__gridTile_35__column__cell.value
          microchart bar #barMicrochart {
            min: 0
            max: 100
            valuePosition: "none"
            colorFormat: SurveyResponseColorScaledMeanScoreFormatter
          }
        }
      }
      column #Dial__gridTile_35__column {
        hide: false
      }
      sort rows #Dial__gridTile_35__sort {
        sortBy: "/Dial__gridTile_35__column"
        sortOrder: "descending"
        takeTop: 20
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: groupOfQuestions
        row: @Dial__gridTile_35__row
        column: @Dial__gridTile_35__column
        cell: @Dial__gridTile_35__column__cell
        sort: @Dial__gridTile_35__sort
        variable: @Dial__gridTile_35__variable
        chartColumn: @Dial__gridTile_35__chartColumn
      }
    }
    size: small
    tile image #imageTile {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20table%20button.png"
      padding: true
      navigateTo: "CX_CS_grid"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_2 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/Trend%20chart%20button.png"
      padding: true
      navigateTo: "CX_CS_trend_line"
      navigateOptions: "same_tab"
    }
    tile image #imageTile_3 {
      value: "/isa/PYAMLMFAKKOYIBEYNHKRJRBIMIEALXOH/KDA%20button.png"
      padding: true
      navigateTo: "CX_CS_KDA_Correlation"
      navigateOptions: "same_tab"
    }
  }
  widget canvas #CX_Comment_divider {
    label: "CX Comment divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "What did members have to say about their overall RX CONCIERGE experience?"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget comments #commentsWidget {
    cardCorners: '20px'
    label: "Please provide any additional comments."
    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: true
      header: surveyDataset_CX:ITLOB
    }
    group question #questionGroup {
      label: "Additional comments"
      filter expression #excludeBlankResponses {
        value: surveyDataset_CX:OA4 != ""
      }
      comment: surveyDataset_CX:OA4
    }
    size: large
    table: surveyDataset_CX:
    cardBackground: #ffffff
    column value #CX_OA1_valueColumn {
      label: "Overall Experience Response"
      value: surveyDataset_CX.response:OA1
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column metric #metricColumn {
      label: "Overall Experience Score"
      value: average(numeric(surveyDataset_CX.response:OA1))
      view: metricView
      target: -1
      align: center
      enableColumnFilter: true
    }
    view metric #metricView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    column value #CX_PlanType_valueColumn {
      label: "Plan Type"
      value: surveyDataset_CX.response:ITPLAN_TY
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #CX_Gender_valueColumn {
      label: "Gender"
      value: surveyDataset_CX.response:ITGENDER
      align: center
      enableColumnFilter: true
      width: "5"
    }
    column value #CX_MemberState_valueColumn {
      label: "Member State"
      value: surveyDataset_CX.response:ITMEMST
      align: center
      enableColumnFilter: true
      width: "5"
    }
  }
  config layout #layoutConfig {
    cardTextColor: "#000000"
    pageBackgroundImage: "None"
  }
  widget canvas #CX_Response_divider {
    label: "CX Survey Response Information divider"
    container: container position {
      width: 1368px
      height: "42px"
      background: #d2ffff
      area #area_4 {
        position: "absolute"
        top: "0px"
        left: "75px"
      }
      area #area_2 {
        position: "absolute"
        top: "-5px"
        left: "13px"
      }
    }
    cardTransparent: true
    tile text #textTile {
      value: "RX CONCIERGE Survey Response Information"
      areaId: "area_4"
      style #style {
        fontSize: 20
        fontFamily: "Arial"
        color: #02253b
        fontWeight: "bold"
      }
    }
    tile image #imageTile {
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/Forsta%20icons/Navy%20icons/Forsta_Icon36.png"
      areaId: "area_2"
      style #style {
        width: "52px"
      }
    }
  }
  widget surveyMetrics #CX_surveyMetricsWidget {
    cardCorners: '20px'
    label: "RX CONCIERGE Survey Metrics"
    mode: "MR"
    scope reportingPeriod #reportingPeriodScope {
      applyTo: "respondent"
    }
    dataSet: surveyDataset_CX
    size: large
  }
  ignoreFilters: fromQuestionFilter_Combo_LOB, fromQuestionFilter_Combo_PLAN, fromQuestionFilter_Combo_CONTRACT, fromQuestionFilter_Combo_GENDER, fromQuestionFilter_Combo_RACE, fromQuestionFilter_Combo_MEMST, fromQuestionFilter_Combo_OA1, fromQuestionFilter_NP_LOB, fromQuestionFilter_NP_PLAN, fromQuestionFilter_NP_CONTRACT, fromQuestionFilter_NP_GENDER, fromQuestionFilter_NP_RACE, fromQuestionFilter_NP_MEMST, fromQuestionFilter_SA_LOB, fromQuestionFilter_SA_PLAN, fromQuestionFilter_SA_CONTRACT, fromQuestionFilter_SA_GENDER, fromQuestionFilter_SA_RACE, fromQuestionFilter_SA_MEMST, fromQuestionFilter_SA_OA1, fromQuestionFilter_AC_LOB, fromQuestionFilter_AC_PLAN, fromQuestionFilter_AC_CONTRACT, fromQuestionFilter_AC_GENDER, fromQuestionFilter_AC_RACE, fromQuestionFilter_AC_MEMST, fromQuestionFilter_AC_OA1, fromQuestionFilter_AC_MA1, fromQuestionFilter_RXCombo_LOB, fromQuestionFilter_RXCombo_PLAN, fromQuestionFilter_RXCombo_CONTRACT, fromQuestionFilter_RXCombo_GENDER, fromQuestionFilter_RXCombo_RACE, fromQuestionFilter_RXCombo_MEMST, fromQuestionFilter_RXCombo_OA1, fromQuestionFilter_RP_LOB, fromQuestionFilter_GP_LOB, fromQuestionFilter_GP_PLAN, fromQuestionFilter_GP_CONTRACT, fromQuestionFilter_GP_GENDER, fromQuestionFilter_GP_RACE, fromQuestionFilter_GP_MEMST, fromQuestionFilter_GP_OA1, fromQuestionFilter_RP_PLAN, fromQuestionFilter_RP_CONTRACT, fromQuestionFilter_RP_GENDER, fromQuestionFilter_RP_RACE, fromQuestionFilter_RP_MEMST, fromQuestionFilter_RP_OA1, fromQuestionFilter_RP_PA4
  hide: true
  modal: false
}




page #CX_OA2_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "RX CONCIERGE NPS"
    series #series {
      value: count(surveyDataset_CX.response:OA2)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: NPSColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_CX:OA2__NPS
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topLeft"
    size: small
    description: "On a scale of 0 to 10, how likely are you to recommend this health plan to a friend or a colleague?"
    layout: "vertical"
  }
  widget headline #CX_Promoters_headlineWidget {
    cardCorners: '20px'
    label: "Promoters"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_CX.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Promoters"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_CX.response:OA2, "10", "9")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Promoters
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Active Promotors are those rating their likelihood to recommend as a 9 or 10"
      size: "small"
    }
  }
  widget headline #CX_Passives_headlineWidget {
    cardCorners: '20px'
    label: "Passives"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_CX.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Passives"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_CX.response:OA2, "8", "7")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Passives
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Passives"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Passives are those rating their likelihood to recommend as a 7 or 8"
      size: "small"
    }
  }
  widget headline #CX_Detractors_headlineWidget {
    cardCorners: '20px'
    label: "Detractors"
    size: small

    tile value #valueTile {
      value: PercentageOfAnswers(surveyDataset_CX.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
    }
    tile text #textTile {
      value: "of members are classified as Detractors"
      fontSize: 18
    }
    tile infographic #infographicTile {
      value: PercentageOfAnswers(surveyDataset_CX.response:OA2, "6", "5", "4", "3", "2", "1", "0")
      valueFormatter: PercentOneDecimalFormatter
      view: iconView_infographicTile
      colorFormatter: colorFormatter_Detractors
    }
    view icon #iconView_infographicTile {
      columns: 10
      rows: 1
      fillDirection: "vertical"
      max: 100
      precision: "exact"
      icon: genderNeutral
    }
    view numeric #numericView_infographicTile {
      max: 100
    }
    infobox #infobox {
      label: "Definition of Active Promotors"
      info: "Likelihood of recommending to friends or colleagues

Scale  0 - 10 (Not at all likely to recommend to Extremely likely to recommend)

Detractors are those rating their likelihood to recommend as 0-6"
      size: "small"
    }
  }
  label: "CX_NPS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #CX_OA1_Stacked_chartWidget {
  widget chart #chartWidget {
    cardCorners: '20px'
    label: "Overall Satisfaction with Rx Concierge"
    series #series {
      value: count(surveyDataset_CX.response:OA1)
      label: "Overall Experience"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_CX:OA1
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    layout: "vertical"
    description: "Overall, I was satisfied with my ability to get appointments for the care I needed."
  }
  label: "CX_OA1 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}





page #CX_OA3_stacked_bar {
  widget chart #CX_OA3_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "RX CONCIERGE - Rating of Health Plan"
    series #series {
      value: count(surveyDataset_CX.response:OA3)
      label: "NPS"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: surveyDataset_CX:OA3
      }
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: large
    description: "Using any number from 0 to 10, where 0 is the worst health plan possible and 10 is the best health plan possible, what number would you use to rate your health plan?"
    layout: "vertical"
  }
  label: "CX_OA3 stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
}




page #CX_CS_stacked_bar {
  label: "CX_CS stacked bar"
  hide: false
  modal: true
  modalSize: "medium"
  widget chart #CX_CS_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rx Concierge"
    series #series {
      value: count(ConRX:value)
      label: "Rx Concierge"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: false
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: ConRX:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
  }
}





page #CX_CS_Components_stacked_bar {
  label: "CX_CS Components stacked bar"
  hide: false
  modal: true
  modalSize: "large"
  widget chart #CX_CS_Components_stacked_bar_chartWidget {
    cardCorners: '20px'
    label: "Rx Concierge Components"
    series #series {
      value: count(ConRX:value)
      label: "Rx Concierge"
      chart bar #barChart {
        mode: "stacked100Percent"
        showBase: false
        showValue: true
        dataLabel: percent
        percentFormat: PercentOneDecimalFormatter
        showBaseInTooltip: true
        maxBarSize: 60
      }
      palette: defaultColorPalette
      format: OneDecimalNumberFormatter

      breakdownBy cut #cutBreakdownby {
        value: ConRX:value
      }
      percentOver: "series"
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: percentScaleNoDecimalDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    legend: "topCenter"
    size: small
    description: ""
    layout: "vertical"
    category cut #cutCategory {
      value: ConRX:field
    }
    chartMargin {
      left: 35
      right: 35
      top: 0
    }
  }
}





page #CX_CS_grid {
  label: "CX_CS grid"
  hide: false
  modal: true
  modalSize: "large"
  widget dataGrid #CX_CS_grid {
    cardCorners: '20px'
    size: large
    column cutByDate #column {
      label: " "
      cell #cell {
        value: average(numeric(ConRX:value))
        view: comparativeStatisticView
        format: OneDecimalNumberFormatter
        showBase: true
      }
      value: surveyDataset_CX:interview_end
      breakdownBy: "calendarMonth"
      showLabel: false
    }
    row cut #row {
      value: ConRX:field
      showLabel: false
      totalLabel: "Rx Concierge"
      label: " "
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: SurveyResponseColorScaledMeanScoreFormatter
      backgroundColorFormatter: SurveyResponseColorPastelBackgroundFormatter
    }
    label: " "
    significanceTesting: true
    confidenceLevels: "95"
    showLegend: false
    fixedHeader: false
  }
}





page #CX_CS_trend_line {
  widget chart #CXtrendchart {
    cardCorners: '20px'
    label: "What are RX MANAGEMENT - Rx Concierge scores over time?"
    chartMargin {
      top: 20
      right: 40
      left: 30
    }
    series #series {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
        showBase: false
      }
      label: "Rx Concierge"
      value: average(numeric(ConRX:value))
      format: OneDecimalNumberFormatter
    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {
      minValue: 0
      maxValue: 100
      format: bigNumberScaleFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
    confidenceLevels: "95"

    selector {
      label: "Trend By"
      option {
        label: "Month"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarMonth

            format: calendarMonthDefaultFormatter
          }
        }
      }
      option {
        label: "Week"
        content {
          category date {
            value: surveyDataset_CX:interview_end
            breakdownBy: calendarWeek
            format: weekFormat
          }
        }
      }
    }
    series #series_2 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Helped save money"
      value: average(numeric(surveyDataset_CX:CX_CS2))
      format: OneDecimalNumberFormatter
    }
    series #series_3 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Made sure taking meds correctly"
      value: average(numeric(surveyDataset_CX:CX_CS3))
      format: OneDecimalNumberFormatter
    }
    series #series_4 {
      chart line #barChart {
        showDotValue: true
        dotSize: 4
        lineType: natural
        lineWidth: 2
      }
      label: "Helped coordinate with provider"
      value: average(numeric(surveyDataset_CX:CX_CS4))
      format: OneDecimalNumberFormatter
    }
    navigateTo: "none"
    description: "RX CONCIERGE - CS Section Scores"
    size: large
    legend: "bottomLeft"
    cardBackground: #ffffff
  }
  label: "CX_CS trend line"
  hide: false
  modal: true
  modalSize: "large"
}





page #CX_CS_KDA_Correlation {
  label: "CX_CS KDA/Correlation"
  hide: false
  modal: true
  modalSize: "large"
  widget keyDrivers #CX_OA2_PA_keyDriversWidget {
    cardCorners: '20px'
    label: "Rx Concierge Key Drivers of NPS (Correlation until enough completes for Regression)"
    size: large
    dependentVariable: surveyDataset_CX:OA2
    independentVariables: surveyDataset_CX:CX_CS2, surveyDataset_CX:CX_CS3, surveyDataset_CX:CX_CS4
    algorithm: correlation
    showOnlySpread: false
    satisfactionLimit: 50.8
    importanceLimit: 0.02
    spreadMode: mean
    cardAlign: center
    cardTransparent: false
    xAxisTitle: "Performance"
    yAxisTitle: "Importance to Members"
    quadrantTitles: "FIX FIRST (Important to Members - Low Scores)", "PROMOTE (Important to Members - High Scores)", "FIX SECOND (Low Importance - Low Scores)", "MAINTAIN(Low Importance - High Scores)"
    cardBackground: #ffffff
  }
  config layout #layoutConfig {
    cardBackgroundColor: ""
  }
}




page #CS {





  label: "CUSTOMER SERVICE"
}





page #COSTS {





  label: "COSTS"
}





page #CAREMGMT {





  label: "RECOMMENDED CARE"
}





page #DISENROLL {





  label: "DISENROLLMENT"
}










config layout #layoutConfig {
  horizontalAlignmentMode: "fullWidth"
  cardTextColor: "#212121"
  pageBackgroundColor: "#ffffff"
}
config breadcrumbs #breadcrumbsConfig {
  combinedText: "Multiple areas of responsibility"
}
