//https://pr.staging.firmglobal.net/apps/editor/191407/summary/
title @externalConfig.reportTitle

// //}





config editor {
  trace: true
}

parameters #externalConfig {
  enduserList: 299
  combinedId: "p620546112173"
  textAnalyticsId: "TextAnalytics_p620546112173_40053"
  reportTitle: "WF test v2"
  usesRespondentFlag: false
  teamIndex1: 4.15
  teamIndex2: 3.8
  leader1: 4
  leader2: 2.5
  numberOfDecimalsForScore: 2
  primaryDimensionId: "engagement"
  filterPanel: layoutArea toolbar {
    filter singleselect #f1 {
      optionsFrom: :EV10040
    }
    filter singleselect #f2 {
      optionsFrom: :EV10013
    }
    filter singleselect #f3 {

      optionsFrom: :EV10022
    }
  }
  demographicsRows: widget dataGrid {
    column {
      hide: true
      cell {
        value: ""
      }
    }
    row cut #EV10013 {
      showLabel: true
      value: :EV10013
      total: first
      collapseMulti: true
    }

    row cut #EV100361 {
      showLabel: true
      value: :EV100361
      total: first
      collapseMulti: true
    }

    row cut #EV10040 {
      showLabel: true
      value: :EV10040
      total: first
      collapseMulti: true
    }

    row cut #EV22864 {
      showLabel: true
      value: :EV22864
      total: first
      collapseMulti: true
    }

    row cut #EV10025 {
      showLabel: true
      value: :EV10025
      total: first
      collapseMulti: true
    }

    row cut #EV10005 {
      showLabel: true
      value: :EV10005
      total: first
      collapseMulti: true
    }

    row cut #EV10020 {
      showLabel: true
      value: :EV10020
      total: first
      collapseMulti: true
    }

    row cut #EV22642 {
      showLabel: true
      value: :EV22642
      total: first
      collapseMulti: true
    }
  }

}

custom properties #cp {
  WFRespondents: count(.respondent:Respondent, .respondent:Respondent = "Yes")
  WFComplete: count(:Respondent, :status = "complete")
  WFResponseRate: @cp.WFComplete / @cp.WFRespondents * 100
}

custom properties #demoPermissions {
  hasSensitive: false
  hasLimited: false
  hasStandard: false
}

reportBase {
  rule nodesKeys {
    reportingHierarchy: unitHierarchy
    values: "Overall"  //root
    //values: "4004454_35278" //leaf
    //values: "4004340_35278" //in beetwen
  }
}

config programNavigation {
  enabled: true
  knowledgeBaseUrl: "https://workforceresources.pressganey.com/"
}

config hub {
  hub: 1628

  referenceData custom #benchmarks {
    table: program_config.benchmark_values:
    selectors: bmValueCode, TrendYear, benchmarkDefinitionID
    array #Per {
      size: 99
    }
  }

  referenceData custom #benchmarksById {
    table: program_config.benchmark_values:
    selectors: bmValueCode, BenchmarkId//, Type
    array #Per {
      size: 99
    }
  }



  reportingHierarchy selfRefLookup #unitHierarchy {
    label: "WF2 to HX newdemo21 - Employee Engagement EV10039"
    source: :EV10039// .respondent:EV10039,  .dg1_questionScore:EV10039 //
    nodeSorting: natural
    showBreadcrumb: true
  }

  dataset custom #project_config {
    publicName: "project_config_" + @externalConfig.combinedId
    defaultTable: report_history //need one to be default
  }


  dataset survey #surveyDataset {
    publicName: @externalConfig.combinedId

    table dimensions = .dg1_dimensions:
    table items = .dg1_questions:
    table benchmarks = project_config.benchmark_list:
    table scaled_items = project_config.scaled_items:
    table dimensionItems = .dg1_dimension_question:
    table rolePermissions = program_config.role_permissions:
    table allPermissions = program_config.allPermissions:
    table widgetConfig = program_config.report_Widgets:
    table reportHistory = project_config.report_history:
    table demo_items = program_config.demo_items:
    table open_items = program_config.open_items:
    table dimension_score = .dg1_dimensionScore:
    table item_score = .dg1_questionScore:
    table dimensionItems = .dg1_dimension_question:




    propagateFilter {
      from: .dimensions:
      to: .dimensionItems:
    }
    propagateFilter {
      from: .dimensionItems:
      to: .items:
    }

    relation oneToMany {
      primaryKey: .scaled_items:itemid
      foreignKey: .items:id
    }

    relation oneToMany {
      primaryKey: .allPermissions:permissionsCode
      foreignKey: .rolePermissions:permissionsCode
    }
    // relation oneToMany {
    //   primaryKey: .reportHistory:prjSurveyPID
    //   foreignKey: :combined_sourceid
    // }
    relation oneToMany {
      primaryKey: .reportHistory:historyTrendOrder
      foreignKey: .item_score:reportHistoryId
    }
    relation oneToMany {
      primaryKey: .reportHistory:historyTrendOrder
      foreignKey: .dimension_score:reportHistoryId
    }
    relation oneToMany {
      primaryKey: .periods:survey
      foreignKey: :combined_sourceid
    }
    relation oneToMany {
      primaryKey: .surveys:code
      foreignKey: :combined_sourceid
    }

    measure custom #dimensionScore {
      value: avg(.dimension_score:dimensionScoreValue)
    }
    measure custom #itemScore {
      value: avg(numeric(.item_score:questionScoreValue))
    }
    // measure custom #itemScoreCount {
    //   value: count(.item_score:)
    // }
    // measure custom #itemScoreSum {
    //   value: sum(numeric(.item_score:questionScoreValue))
    // }

    variable numeric #forDimension {
      table: :
      value: avg(.dimension_score:dimensionScoreValue, .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId, :)
    }


   //TODO: can we get rid of this hardcoding?
    recoding ranges #LeaderIndexGroup {
      intervals: leftopen
      mapping {
        to: "Low"
        from: "..3"
      }
      mapping {
        to: "Moderate"
        from: "3..4"
      }
      mapping {
        to: "High"
        from: "4.."
      }


    }


  }

  dataset textAnalytics #textAnalyticsDataset {
    publicName: @externalConfig.textAnalyticsId
    table responses = surveyDataset.response:
  }
  dataSet: surveyDataset



  //Selector content for response rate page
  dataTable #dtResponseRateItems {
    dataGrid #dgresponseRateItems {
      size: large
      row #rritems {
        row #orgunithier {
          cell custom {
            expression #id {
              value: "EV10039"
            }
            expression #label {
              value: "Organization hierarchy - Hierarchy"
            }
            expression #rows {
              value: "hier"
            }
            expression #cols {
              value: "invited, responded, rate"
            }
            formatString: "{id} {label}"
          }
        }
        row #orgunit {
          cell custom {
            expression #id {
              value: "EV10039"
            }
            expression #label {
              value: "Organization hierarchy - Flat"
            }
            expression #rows {
              value: "units"
            }
            expression #cols {
              value: "invited, responded, rate, rollup" //"rollup"
            }
            formatString: "{id} {label}"
          }
        }
        //TODO: Only list demographics user have access to!   
        row list #demos {
          total: none
          table: .demo_items:
          value: ""
          filter expression {
            value: .demo_items:cmbdSurveyPID = @externalConfig.combinedId
          }
          cell custom {
            expression #id {
              value: .demo_items:itemID
            }
            expression #label {
              value: .demo_items:itemLabel
            }
            expression #rows {
              value: "cut"
            }
            expression #cols {
              value: "invited, responded, rate"
            }
            formatString: "{id} {label}"
          }
        }
      }
      column #main {

      }
    }
    map #forSelect2 {
      from: "rritems"
      to: item {
        label: this.main.label
        value:  {
          id: this.main.id
          col: studio.expressionFromCdl(this.main.cols)
          row: this.main.rows
        }
      }
    }
  }

  //Calculating available rollup modes depending on where in the hierarchy user is
  dataTable #dtModes {
    dataGrid #dgModes {
      removeEmptyRows: true
      row #nodes {
        //hide: true
        cell {
          value: IIF(count(unitHierarchy:) != countIf(IsLeaf(unitHierarchy:^hierarchy)), "PARENT", "LEAF")
        }
      }

      row #variants {
        row #v1 {
          cell custom {
            formula #label {
              value: IIF([row = /nodes] = "PARENT", "My Team View")
            }
            formula #mode {
              value: IIF([row = /nodes] = "PARENT", "rollup")
            }
            formula #gridMode {
              value: IIF([row = /nodes] = "PARENT", "rollup")
            }
            formatString: "{label} {mode} {gridMode}"
          }
        }
        row #v2 {
          cell custom {
            formula #label {
              value: IIF([row = /nodes] = "PARENT", "Direct Reports")
            }
            formula #mode {
              value: IIF([row = /nodes] = "PARENT", "direct")
            }
            formula #gridMode {
              value: IIF([row = /nodes] = "PARENT", "mixed")
            }
            formatString: "{label} {mode} {gridMode}"
          }
        }
        row #v3 {
          cell custom {
            formula #label {
              value: IIF([row = /nodes] = "LEAF", "My Team (as Direct)")
            }
            formula #mode {
              value: IIF([row = /nodes] = "LEAF", "direct")
            }
            formula #gridMode {
              value: IIF([row = /nodes] = "LEAF", "mixed")
            }
            formatString: "{label} {mode} {gridMode}"
          }
        }
      }
      column #status {
      }
    }
    map #forSelect {
      from: "variants"
      to: item {
        label: this.status.label
        value:  {
          mode: this.status.mode
          gridMode: this.status.gridMode
        }
      }
    }
  }

  dataTable #dtOpenItems {
    dataGrid #dgOpenItems {
      filter expression {
        value: .open_items:cmbdSurveyPID = @externalConfig.combinedId
      }
      row list #open {
        total: none
        table: .open_items:
        value: ""
      }
      column #main {
        cell custom {
          expression #id {
            value: .open_items:itemID
          }
          expression #label {
            value: .open_items:itemLabel
          }
          formatString: "{id} {label}"
        }
      }
    }
    map #forSelect {
      from: "open"
      to: item {
        label: this.main.label
        value: this.main.id
      }
    }
  }

  dataTable #dtEngagementSummary {
    dataGrid #dgEngagementSummary {
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      // filter expression {
      //   value: .reportHistory:cmbdSurveyPID = @externalConfig.combinedId
      // }

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }

      row #engagement {
        filter expression {
          value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
        }
      }

      column cut #history {
        scope filter {
          name: period
          value: currentAndPrevious
        }
        value: .reportHistory:historyTypeCode
        total: none

        cell custom {
          expression #score {
            value: :dimensionScore()
            //formatter: numberFormatter_5
          }
          statistic mean #sig {
            testingType: T
            argument: .dimension_score:dimensionScoreValue
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diff}"
        }
      }
      column #main {
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
          }
          formula #sig {
            value: sig[column = /history.current]
          }
          formula #asteric {
            value: IIF(sig[] != 0, "*", " ")
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #sigInfo {
            value: IIF(sig[] != 0, "change is statistically significant", "change is not statistically significant")
          }
          formatString: "{current} ({change}) [{sig}]"
        }
      }

      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarksById
            mapping value {
              value: @externalConfig.primaryDimensionId
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.idInt
              selector: BenchmarkId
            }
            value: :dimensionScore()
            formatter: rankFormatter
          }
          formatString: "{rank}"
        }
      }
      column #microchart {
        cell microchart {
          value: count(.dimension_score:)
          breakdownBy cut {
            value: .dimension_score:engagementFourPoint
          }
          microchart pie {
          }
        }
      }
    }

    map #m {
      from: engagement
    }
  }


  dataTable #rolePermissions {
    dataGrid {
      filter expression {
        value: .rolePermissions:cmbdSurveyPID = @externalConfig.combinedId AND .rolePermissions:roleCode = @userRole.selected
      }

      column #permission {
        cell {
          value: .allPermissions:permissionsCode
        }
      }
      column #permissionCount {
        cell {
          value: count(.rolePermissions:permissionsCode)
        }
      }
      column #isHidden {
        cell {
          value: count(.rolePermissions:permissionsCode) = 0
        }
      }
      row list #permissions {
        table: .allPermissions:
        value: .allPermissions:permissionsCode

      }


    //  map #forSelect {
    //   from: "permission"
    //   to: {
    //     permission: this.permission.value
    //   }
    // }
    }
    map #permissionLookup {
      from: "permissions"
      to:  {
        permission: this.permissionCount.value
        isHidden: this.isHidden.value
      }
      toRecord byKey {
        key: this.permission.value
      }
    }

  }

  dataTable #widgetConfig {
    dataGrid {
      label: "Data Grid"
      size: "large"
      filter expression {
        value: .rolePermissions:cmbdSurveyPID = @externalConfig.combinedId
      }
      column #widgetCode {
        cell {
          value: .widgetConfig:widgetCode
        }
      }
      column #widgetLabel {
        cell {
          value: .widgetConfig:widgetLabel
        }
      }
      column #widgetDescription {
        cell {
          value: .widgetConfig:widgetDescription
        }
      }
      column #widgetInfoText {
        cell {
          value: .widgetConfig:widgetInfoText
        }
      }
      row list #widgetCodes {
        table: .widgetConfig:
        value: .widgetConfig:widgetCode
      }
    }
    map #lookup {
      from: "widgetCodes"
      to:  {
        label: this.widgetLabel.value
        description: this.widgetDescription.value
        infoText: this.widgetInfoText.value
      }
      toRecord byKey {
        key: this.widgetCode.value
      }
    }
  }

  //dataTable getting list of dimensions from table .dimensions: to fill in selectors, including what is default
  dataTable #dtDimensions {
    dataGrid #dgDimensions {
      row list #dimensions {
        total: none
        table: .dimensions:
        value: ""
        sortBy: "/_label"
        sortOrder: ascending
      }

      column #results {
        cell custom {
          expression #label {
            value: .dimensions:id //[column = /_label]
          }
          expression #type {
            value: "leader" //.dimensions:typeMG
          }
          expression #id {
            value: toText(.dimensions:id)
          }
          expression #isDefault {
            value: .dimensions:isPrimary
          }
          formula #points {
            value: IIF(type[] = "Engagement", "fourPoint", "threePoint")
          }
          formatString: "{label} | {type} | {id} | {isDefault}"
        }
      }
    }
    map #forSelect {
      from: "dimensions"
      to: item {
        label: this.results.id
        value:  {
          id: this.results.id
          type: this.results.type
          isDefault: this.results.isDefault
          points: this.results.points
        }
      }
    }
    map #forSelect2 {
      from: "dimensions"
      to: item {
        label: this.results.label
        value: this.results.id
        isDefault: this.results.isDefault
      }
    }
  }
  dataTable #dtItems {
    dataGrid #dgItems {
      row list #items {
        total: none
        table: .items:
        value: ""
        sortBy: "/num"
        sortOrder: ascending
      }
      column #num {
        hide: true
        cell {
          value: .items:sequenceId
          extraValue: toText(.items:sequenceId)
        }
      }
      column #results {
        cell custom {
          expression #label {
            value: .items:label
          }
          formula #fullLabel {
            value: extraValue[column = /num] + ". " + label[]
          }
          expression #id {
            value: toText(.items:id)
          }
          formatString: ""
        }
      }
    }
    map #forSelect {
      from: "items"
      to: item {
        label: this.results.fullLabel
        value: this.results.id

      }
    }
  }
  dataTable #dtSurveys {
    dataGrid #dgSurveys {
      row list #surveys {
        filter expression {
          value: .reportHistory:historyTrendOrder != 1

        }
        total: none
        table: .reportHistory:
        value: ""
      }
      column #col {
        cell custom {
          expression #id {
            value: .reportHistory:historyTrendOrder
          }
          expression #label {
            value: .reportHistory:historyLabel
          }
          expression #code {
            value: .reportHistory:prjSurveyPID
          }
          expression #isDefault {
            value: .reportHistory:historyTrendOrder = 2
          }
          expression #trendOrder {
            value: toText(.reportHistory:historyTrendOrder)
          }
          formatString: ""
        }
      }
    }
    map #forSelect {
      from: surveys
      to: item {
        label: this.col.label
        value: this.col.id
        isDefault: this.col.isDefault
        trendOrder: this.col.trendOrder
      }
    }
  }
  dataTable #dtBenchmarks {
    dataGrid {
      row list #benchmarks {
        total: none
        table: .benchmarks:
        value: ""
        sortBy: "/order"
        sortOrder: ascending
      }
      column #order {
        hide: true
        cell {
          value: .benchmarks:benchmarkOrder
        }
      }
      column #results {
        cell custom {
          expression #label {
            value: .benchmarks:benchmarkName
          }
          expression #id {
            value: .benchmarks:BenchmarkID
          }
          expression #idText {
            value: toText(.benchmarks:BenchmarkID)
          }

          expression #definitionId {
            value: .benchmarks:BenchmarkDefinitionID
          }
          expression #definitionName {
            value: .benchmarks:BenchmarkDefinitionName
          }
          expression #periodId {
            value: .benchmarks:TrendYear
          }
          expression #order {
            value: toText(.benchmarks:id)
          }
          formatString: "{label} {definitionId} {isDefault}"
        }
      }
    }
    map #forSelect {
      from: "benchmarks"
      to: item {
        label: this.results.label
        value: this.results.id
        idText: this.results.idText
  //      order: this.results.order
      }
    }
  }


}

config queryOptions {
  // added automatically during report creation
  boolNullsAsFalse: false
  explicitLevelAggregation: false
}

layoutArea toolbar @externalConfig.filterPanel { //
  useDynamicFilters: true

  filter singleselect #isRespondentFilter {
    label: "IsRespondentFilter"
    hide: true
    option checkbox {
      label: "Respondent=YES"
      value: :respondent = 'YES'
      selected: @externalConfig.usesRespondentFlag

    }
    option checkbox {
      label: "No Respondent Filter"
      value: true
      selected: @externalConfig.usesRespondentFlag = false
    }

  }
  filter reportingHierarchy #unitHierarchyFilter {
    reportingHierarchy: unitHierarchy
    label: "Unit Hierarchy"
  }
  filter singleselect #cur {
    //label: "Current"
    scope {
      name: period
    }
    hide: true
    option radio #current {
      //label: "current"
      //value: .reportHistory:historyTypeCode = "current"
      value: .reportHistory:historyTrendOrder = 1
      selected: true
    }
  }
  filter singleselect #curAndPrev {
    scope {
      name: period
      value: currentAndPrevious
    }
    hide: true
    option radio #currentAndPrevious {
      //value: .reportHistory:historyTypeCode = "current" OR .reportHistory:historyTypeCode = "primary"
      value: .reportHistory:historyTrendOrder = 1 OR .reportHistory:historyTrendOrder = 2
      selected: true
    }
  }
  filter singleselect #prev {
    scope {
      name: period
      value: previous
    }
    hide: true
    option radio #previous {
      value: .reportHistory:historyTypeCode = "primary"
      selected: true
    }
  }

  widget toolbarWidget {
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      mode: @rollupMode.selected.mode
    }
    tile custom {
      expression #first {
        value: @cp.WFComplete
        formatter: bigNumberFormatter
      }
      expression #second {
        value: @cp.WFComplete / COUNT(:responseid) * 100
        formatter: percentNoDecimal
      }
      fontSize: 16
      formatString: "{first} Responses ({second})"
    }
    select #rollupMode {
      //label: "Rollup mode e"
      options: @dtModes.forSelect.data
    }
  }
}

config style #styleConfig {
  theme: "modern"
}

config report {
  formatter number #scoreFormatter {
    decimalSeparator: "."
    numberDecimals: @externalConfig.numberOfDecimalsForScore
    integerSeparator: ","
    emptyValue: "-"
    keepTrailingZeros: true
  }
  formatter number #diffFormatter {
    decimalSeparator: "."
    numberDecimals: @externalConfig.numberOfDecimalsForScore
    integerSeparator: " "
  }
  formatter number #rankFormatter {
    ordinal: true
    emptyValue: "-"
    integerSeparator: ","
    numberDecimals: 0
  }

  formatter color #taSentimentColorFormatter {
    label: "Red Amber Green (Sentiment)"
    thresholds: #1DA583 > 0.25, #E79F0D >= -0.25, #d02525 >= -5
  }
  formatter color #taSentimentDefaultBackgroundColorFormatter {
    label: "TA Sentiment Background Color Numeric"
    thresholds: #D3EFDA > 0.25, #FFFFE0 >= -0.25, #F7D4D4 >= -5
    defaultValue: #FFFFE0
  }
  formatter color #positiveColorDefaultFormatter {
    label: "Positive"
    thresholds: #1DA583 > 0
  }
  formatter color #neutralColorDefaultFormatter {
    label: "Neutral"
    thresholds: #E79F0D > 0
  }
  formatter color #negativeColorDefaultFormatter {
    label: "Negative"
    thresholds: #d02525 > 0
  }
  formatter color #sentimentindicatortextValue {
    thresholds: Positive > 0, Neutral = 0, Negative < 0
  }
  formatter color #sentimentindicator {
    thresholds: #1DA583 > 0, #E79F0D = 0, #d02525 < 0
    defaultValue: transparent
  }
  formatter color #sentimentindicatortext {
    thresholds: #FFFFFF > 0, #333333 = 0, #FFFFFF < 0
  }

  formatter date #dayformatter {
    formatString: "ddd, MMM DD"
  }
  formatter number #bigNumberFormatter {
    label: "integerFormatter"
    numberDecimals: 0
    prefix: ""
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: false
    ordinal: false
  }
  formatter number #floatDefaultFormatter {
    label: "two_decimalsFormatter"
    numberDecimals: 2
    prefix: ""
    postfix: ""
    decimalSeparator: "."
    integerSeparator: ","
    shortForm: false
    keepTrailingZeros: true
    ordinal: false
  }
  palette answerList #LIpalette {
    hint visualDesigner #visualDesignerHint {
      type: "answerListPalette"
      value: .response:LeaderIndexGroup
    }
    item #item {
      code: "High"
      color: #1FA583
    }
    item #item_2 {
      code: "Moderate"
      color: #E79F0B
    }
    item #item_3 {
      code: "Low"
      color: #D02525
    }
    label: "Leader Index Palette ee"
  }
  palette answerList #engaged { //colors4 CNJ 
    item {
      code: "4"//"Disengaged"
      color: #D75D38
    }
    item {
      code: "1"//"Highly Engaged"
      color: #027580
    }
    item {
      code: "2"//"Engaged"
      color: #1FA583
    }
    item {
      code: "3"//"Neutral"
      color: #E79F0B
    }

  }
  palette answerList #favorable { //colors3 CNJ
    item {
      code: "3"//"Unfavorable"
      color: #D02525
    }
    item {
      code: "1"//"Favorable"
      color: #1FA583
    }
    item {
      code: "2"//"Neutral"
      color: #E79F0B
    }

  }
  palette #ragPalette {
    colors: "#1DA583","#E79F0D","#d02525"
    label: "Red Amber Green (Palette)"
  }
}

config pdfExport {
  pageSize: A4, A3, Letter
  pageOrientation: portrait, landscape
  pageScaling: fitToWidth
  exportMode: htmlToPdf
  version: 2
  allowFileNaming: true
  pageMargins: 0.4
}

config mobile {
  showShareButton: true
}

page #Page1 {
  hide: true
  label: "Settings"
  widget headline {
    label: "Hardcoded selectors - USE THEM"
    size: large
    tile text #textTile_2 {
      value: "What is selected here is applied to all pages"
    }
    select #userRole {
      label: "Role"
      options: item { label: "pgfAdmin" value: "pgfAdmin"},
      item {label: "DefaultManager" value: "DefaultManager"},
      item {label: "defaultViewAll" value: "defaultViewAll"},
	    item {label: "defaultLeader" value: "defaultLeader"},
	    item {label: "hr" value: "hr"}
      defaultOption: "defaultViewAll"
    }
    //This one is moved to toolbar
    // select #rollupMode {
    //   label: "Rollup mode"
    //   options: item { label: "My team view" value: {mode: rollup gridMode: rollup}},
    //   item {label: "Direct view" value: {mode: direct gridMode: mixed}},
    //   item {label: "My team view as direct" value: {mode: direct gridMode: direct}}
    // }
    select #defaultBenchmmark {
      label: "Default benchmark"
      options: item { label: "Nat'l Healthcare Avg (Employee) 2023" value: {idText: "3871" idInt: 3871 definitionId: 2 definitionName: "Nat'l Healthcare Avg" periodId: 2023 } },
      item { label: "Nat'l Academic Healthcare Avg 2023" value: {idText: "3879" idInt: 3879 definitionId: 3 definitionName: "Nat'l Academic Avg" periodId: 2023 } },
      item { label: "Nat'l Healthcare Avg (Employee) 2020" value: {idText: "3430" idInt: 3430 definitionId: 2 definitionName: "Nat'l Healthcare Avg" periodId: 2020 } },
      item { label: "Nat'l Healthcare Avg (Employee) 2019" value: {idText: "3095" idInt: 3095 definitionId: 2 definitionName: "Nat'l Healthcare Avg" periodId: 2019 } }
    }
    select #surveyToCompareWith {
      //MG if no previouis survey use the current but hide columns
      label: "Survey to compare with"
      options: item { label: "Employee Engagement 2020" value: {id: 2 code: p217979574846 } },
      item { label: "Employee Engagement 2021 - DO NOT SELECT" value: {id: 1 code: p494984785246 } }
    }
    select #suppressionThreshold {
      label: "min Sample Size"
      options: item{ label: "1" value: 1}, 
      item{ label: "10" value: 10},
      item{ label: "25" value: 25},
      item{ label: "50" value: 50},
      item{ label: "100" value: 100}
    }
  }

  //   widget headline #headlineWidget_3 {
  //   label: "That are properly filled in selectors - DON'T USE THEM - waiting for #3"
  //   size: large
  //   tile text {
  //     value: "What is selected here is applied to all pages"
  //   }
  //   select #rollupMode1 {
  //     label: "Rollup mode"
  //     options: @dtModes.forSelect.data
  //   }
  //   select #defaultBenchmmark1 {
  //     label: "Default benchmark"
  //     options: @dtBenchmarks.forSelect.data
  //     defaultOption: true
  //     compareBy: this.value.isDefault
  //   }
  //   select #surveyToCompareWith1 {
  //     label: "Survey to compare with"
  //     options: @dtSurveys.forSelect.data
  //   }
  //   select #suppressionThreshold1 {
  //     label: "min Sample Size"
  //     options: item{ label: "1" value: 1}, 
  //     item{ label: "10" value: 10},
  //     item{ label: "25" value: 25},
  //     item{ label: "50" value: 50},
  //     item{ label: "100" value: 100}
  //   }
  // }

  widget markdown #cl {
    size: large
    label: "Change log - create new document revision before making major changes"
    markdown: "    * FW 2/2: Remove old, deprected Items, fixed scope for widget toolbarWidget
    * 2/1 DHE: Added CA Modal, Split EI and Leader Widgets (Summary, Overall, DR)
    * 2/1 FW: Set default role to defaultViewAll
    * 1/31 DHE: Added the Overall Page
    * 1/31 FW: Exclude items from key driver
    * 1/30 FW: Using new project specific tables for report_history and benchmark_list
    * 1/29 DHE: Edited Direct report Engagement trend to show.
    * 1/29 DHE: Edited summary arrows.
    * 1/29 DHE: Edited Demo Performance widgets.
    * 1/29 DHE: Added Direct Report Summary widgets
    * 1/29 FW: Added global filter for report_history on cmbdSurveyPID
    * 1/28 DHE: Added Palette for CA. **Note this has an issue where one of the colors is not coming through**
    * 1/28 CMB: Updated Leader Index, references.
    * 1/28 JFA: change supress rule expression - reportHistory.id = 1001 TODO: Needs to fix logic
    * 1/26 DHE: Updated Leader Index with score. **NOTE: Still needs calculations for the High/Moderate/Low text underneath** 
    * 1/26 CNJ: legend on 5 donuts  
    * 1/26 CNJ: 5 donuts in a row. see //CNJ126 tileset 
    * 1/26 DylanE: Updated Key Drivers Mean score to include arrow and Sig. Added Top Performers Widget.
    * 1/26 DylanE: Change Key Drivers Format to remove decimals
    * 1/26 CNJ: Changes on Engagement widget; replaced container, added legend , modified chart
    * 1/26 CNJ: - changes across summary page to keep one legend type (diamond, it was the one that got better aligned as a legend on engagement) see “CNJ126 legend”. Consider changing legend all across for consistency
    * 1/26 CNJ: cleaned up code
    * 1/26 CNJ: prettified arrows, and adjusted text in donuts - CNJ126 arrows
    * 1/25 Carolyn: Updated suppression messages.  minor edits.
    * 1/25 DylanE: Changed Hovers for summary widgets, added sig color to Eng for lrg groups.
    * 1/25 DylanE: Updated overall tool bar responses formatting and added too few suppression to summary widgets
    * 1/24 DylanE: Updated Hover functionality, Sig Score Color, Colors to charts
    * 1/24 DylanE: Updated Additional Experience Dimensions Widget and Updated all summary widgets to display based on ʺMy Team Viewʺ vs ʺDirect Reportʺ
    * 1/24 FrankW: added support for Respondent=YES filter via CDL parameters
    * 1/23 DylanE: Updated Summary Widgets ( Response Rate, Engagement, Leader Index,Engagement Largest groups, Engagement Trend, Key Drivers of Engagement) 
    * 01/20 FrankW: Fixed demographic selector on ResponseRate
     
    
      Leade"

  }

  widget markdown #todo {
    size: large
    label: "TODO"
    markdown: "Frank / Mikhail
- fix trend chart on Summary page -- only showing current values.
- Selectors for Item Details
- Selectors for Org Details and Demographic Details
- setting for Overall Organization page (not yet added) so that the results always reflect top full organization results, 

- Find a way to only show this settings page for professional users (I will hide page for the Monday demo)
- Exclude items from key drivers calculation - FrankW -- (note, I manually excluded these in the CDL, but the calculations need to be updated to only use the correct items from the custom data table.)
- ~~Key Demographics calculation~~
-~~ Update widget table to reference this report.  I added all of the widgets to the table -- validate with Joffe~~
- How should we display hovers of suggested actions

- ~~Address duplicate combined surveys and impact into individual reports (doubles responses for current survey)~~
- Roles and levels in the hierarchy - what to do when navigating to lowest level (but not assigned to that level), switch to DR only?
-Thomas - nesting in the crosstab
- Verify how to set up the heatmaps in crosstab and/or details pages and associate to views in the selectors?
- Questions for the suppression rules, specifically when the too few is for individual items / rows and not for the entire team.
- deploy to production / enable toggles in WF Company on HX

Outstanding layout / look & feel
~~-Summary - Spacing Engagement widget, display legend CNJ~~
~~-Cleaner arrows, with more space between mean score and arrow in tables.  Arrow needs to continue to support colors for significance.~~
~~-JV's feedback for the Largest Group widget (five donuts in a row) -   display legend~~
-~~Add Leader Index mean score and category (High, Medium, Low) to the Leader Index widget.  I added three areas, but formatting is still needed.~~
~~- On Key Drivers, correct hover (remove decimals)~~
~~- Key Drivers, add sig arrow to Mean score~~
- Incorporate selector example from 191198 on Item details
- Fix comment analytics legend, switch to 3 column 
- Update description fields
-Additional layout and alignment
-Refresh snapshot with updated widgets
- duplicate for DR and overall
- Key Demographics, Team Index, Alignment/Engagement combo, eNPS, 

Fix
- Trend chart not showing values
~~- Dylan - add Top Performers once we verify we should add widget references for the template~~







Calculations
-Exclude items from key drivers
-Key Demographics
~~-Top Performers - DHE: Waiting on the label, info, and description to be put in.~~

Summary
- Megan - All widgets, address spacing between Title and Description (increase font??)

Questions/Assistance / Status

1. Selectors (Mikhail)
--noticed in the modal that dimension are displaying the code, not the label
--fixed in 191198
2. Exclude items from key driver analysis based on configuration (Frank)
3. Key demographic calculation (Frank)
~~4. How to address suppression issues / message~~
5. Click throughs from Summary using the selectors on item details, work unit, demographics - ensure correct dimensions selected
6. Display two horizontal bar graphs in single widget instead of vertical bar graphs - or do we have to have two separate widgets?
~~7. Cannot get the legend to display for donut now that it is a micro chart~~
~~8. Number formatter not working on toolbar # of responses~~
9. Is there any way to update the content within chart hovers? e.g. percentage displays, but tag is number of responses
~~10. How do we get the headers to display at the top of each column within tables?~~ 
11. What options do we have to better format the list tables?
12. Update arrows for statistical significance -- bigger.  Can we have more space between mean score and arrows?
~~13. Update the number formatters in the chart hover overs~~
14. How should suggested action hovers be set up for the individual items?
~~16. Dylan - need to review the hover over changes, getting mean scores not calculating.  I have not merged my updates.~~
17. How do we keep Overall Organization page to always reflect top level of hierarchy?
~~18. Dylan - are you good with how to display different widgets when Direct Reports selected?  and vice versa with My Team View?~~
19.  What is the format we need to apply for the roles?


Meeting requested with JV
~~- Add correct suppression messages , hide items, charts, comparisons~~
~~- Add colors to statistical significance~~
- legends
- bottom padding
~~- add Top Performers (copy Key Drivers, change calc)~~
- add Key Demographics
- add Team Index (copy Leader Index)
- create Direct Reports versions for widgets, associate to drop down
- create Overall Organization version for widgets
- add click throughs (after selectors and modals added to Items, Work Units, and Demographics)

Engagement Widget
~~- Update donut with correct colors~~
- Add legend
- Shift chart and table (space from the center)
- Update hover format / content for table

Trend
-Display only My Team if at top level

Leader Index
~~- Add score and category~~
~~- Shift to three areas~~

Largest Groups
~~- Apply correct colors~~
~~- add ʺPercentileʺ after percentile~~
~~- Responses, not Respondents~~

Key Drivers
- Apply correct colors to response distribution
~~- Update hover to include thousands comma~~
- Add hover to item with the suggested action

Related HX Dimensions
- Hide column with TI-2
- align values under headers

Items
-  Set selectors (view, display, dimensions)
- Modal
- Responds to Direct Reports
- Suppression messages

Work Unit
-  Set selectors (view, display, dimensions)
- Modal
- Responds to Direct Reports
- Suppression messages"

  }



  //dataTable #dtBenchmarks {
  // widget dataGrid #dgBenchmarks {
  //   row list #benchmarks {
  //     total: none
  //     table: .benchmarks:
  //     value: ""
  //     sortBy: "/published"
  //     sortOrder: descending
  //   }
  //   column #published {
  //     hide: true
  //     cell {
  //       value: .benchmarks:benchmarkDate
  //     }
  //   }
  //   column #results {
  //     cell custom {
  //       expression #label {
  //         value: .benchmarks:benchmarkName
  //       }
  //         // expression #id {
  //         //   //MG it is "single" in benchmark table but int in benchmarkValues table
  //         //   value: toText(.benchmarks:BenchmarkID)
  //         //   //value: .benchmarks:BenchmarkID
  //         // }
  //       expression #idInt {
  //         value: .benchmarks:BenchmarkID
  //       }
  //       expression #definitionId {
  //         value: .benchmarks:BenchmarkDefinitionID
  //       }
  //       expression #definitionName {
  //         value: .benchmarks:BenchmarkDefinitionName
  //       }
  //       expression #periodId {
  //         value: .benchmarks:TrendYear
  //       }
  //       expression #isDefault {
  //         value: .benchmarks:benchmarkIsPrimary
  //       }
  //       formatString: "{label} {idInt} {definitionId} {isDefault}"
  //     }
  //   }
  // }
  // map #forSelect {
  //   from: "benchmarks"
  //   to: item {
  //     label: this.results.label
  //     value:  {
  // //        id: this.results.id
  //       isDefault: this.results.isDefault
  //       idInt: this.results.idInt
  //       definitionId: this.results.definitionId
  //       definitionName: this.results.definitionName
  //       periodId: this.results.periodId
  //     }
  //   }
  // }
  //}


}
page #summary {

  label: "Summary"
  scope reportingHierarchy {
    reportingHierarchy: unitHierarchy
    mode: @rollupMode.selected.mode
  }
  dataTable #dtEngagementNodes {
    dataGrid #dgEngagementNodesTMP {

      scope filter {
        name: period
        value: currentAndPrevious
      }

      size: large
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }
      filter expression {
        value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
      }

      row list #nodes {
        total: none
        table: unitHierarchy:
        value: ""//unitHierarchy:language_text
        // takeTop: 5
        // sortBy: "/base"//count(:, .surveys:id = 1)
        take: 5
        sortBy: count(:, .reportHistory:historyTypeCode = "current")
        sortOrder: descending
      }

      column #nodeLabel {
        cell {
          value: unitHierarchy:language_text
        }
      }
      column #base {
        cell {
          value: count(:, .reportHistory:historyTypeCode = "current")
        }
      }
      column cut #history {
        // scope filter {
        //   name: period
        //   value: currentAndPrevious
        // }
        value: .reportHistory:historyTrendOrder
        total: none

        cell custom {
          expression #score {
            value: :dimensionScore()
          }
          statistic mean #sig {
            testingType: T
            argument: .dimension_score:dimensionScoreValue
            compare: next
          }

          formatString: "{score} [{sig}]"
        }
      }
      column #main { //This is where Engagement For your largest Groups is obtained from
        label: main
        cell custom {
          formula #score {
            value: score[column = /history.1]
          }
          formula #change {
            value: score[column = /history.1] - score[column = /history.2]
          }
          formula #sig {
            value: sig[column = /history.1]
          }
          formula #asteric {
            value: IIF(sig[] != 0, "*", " ")
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #historyMean {
            value: score[column = /history.2]
          }
          formula #sigInfo {
            value: IIF(sig[] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.1] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.1] != 0, "#d02625", "Black"), "Black"))
          }
          formatString: "{score} ({change}) [{sig}]"
        }
      }

      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarksById
            mapping value {
              value: @externalConfig.primaryDimensionId
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.idInt
              selector: BenchmarkId
            }
            value: :dimensionScore()
            formatter: rankFormatter
          }
          formatString: "{rank}"
        }
      }
      column #microchart {
        cell microchart {
          value: count(.dimension_score:)
          breakdownBy cut {
            value: .dimension_score:engagementFourPoint
          }
          microchart pie {
          }
        }
      }
    }
    map #m {
      from: nodes
    }
  }

  // widget toolbarWidget #page1Toolbar {
  //   size: large

  //   tile custom {
  //     expression #first2 {
  //       value: @cp.WFComplete
  //     // formatter: noDecimalsUS
  //     }
  //     expression #second2 {
  //       value: @cp.WFComplete / @cp.WFRespondents * 100
  //       formatter: percentNoDecimal
  //     }
  //     fontSize: 16
  //     formatString: "Select Benchmark"
  //   }
  //   // select #rollupMode2 {
  //   //   // label: "Rollup mode"
  //   //   options: item { label: "My team view" value: {mode: rollup gridMode: rollup}},
  //   //   item {label: "Direct view" value: {mode: direct gridMode: mixed}},
  //   //   item {label: "My team view as direct" value: {mode: direct gridMode: direct}}
  //   // }
  //   select #defaultBenchmmarkSummary {
  //     // label: "Benchmark"
  //     options: item { label: "Nat'l Healthcare Avg (Employee) 2021" value: {idInt: 3871 definitionId: 2 definitionName: "Nat'l Healthcare Avg" periodId: 2021 } },
  //     //updated the label for 3430 just for the purposes of the demo.  
  //     item { label: "Nat'l Academic Avg 2021" value: {idInt: 3430 definitionId: 2 definitionName: "Nat'l Healthcare Avg" periodId: 2020 } }
  //     //item { label: "Nat'l Healthcare Avg (Employee) 2019" value: {idInt: 3095 definitionId: 2 definitionName: "Nat'l Healthcare Avg" periodId: 2019 } }
  //   }

  //   // select #defaultBenchmmarkNew {
  //   //   label: "Default benchmark"
  //   //   options: @dtBenchmarks.forSelect.data
  //   //   defaultOption: true
  //   //   compareBy: this.value.isDefault
  //   // }

  //   // select #MyTeamViewSelector {
  //   //   background: transparent
  //   //   options: item {
  //   //       label: "My Team View"
  //   //       value: false
  //   //    },
  //   //   item {
  //   //       label: "My Direct Reports"
  //   //       value: true
  //   //  // },
  //   //  //  item {
  //   //  //     label: "Overall Organization View"
  //   //    //   value: true
  //   //   }
  //   // }

  // }



  widget headline #summaryMTVResponseRate {
    label: @widgetConfig.lookup.data.summaryMTVResponseRate.label
    description: @widgetConfig.lookup.data.summaryMTVResponseRate.description
    size: large
    hide: @rollupMode.selected.mode != "rollup"

    // Do not need to hide values on response rate widget
    // suppressRule {
    //   criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
    //   label: "Too few responses" //what to display
    // }
    // hide: @rollupMode.Selected.value

    toolbar { //start toolbar
      button #infobox {
        action showInfobox {
          info: @widgetConfig.lookup.data.summaryMTVResponseRate.infoText
          label: @widgetConfig.lookup.data.summaryMTVResponseRate.label
          size: large
        }
      }
      button #export {
        action export {
          format: png
        }
      }
      button #navigate {
        action navigate {
          navigateTo: response_rates
        }
      }
    } //end toolbar
    container: container flex {
      flexDirection: row
      flexWrap: wrap

      area #area_one_space {
        width: '7%'
        display: block
      }
      area #area_one {
        width: '9%'
        display: block
        verticalAlign: "center"
      }
      area #area_two {
        width: '13%'
        display: block
      }
      area #area_three_space {
        width: '12%'
        display: block
      }
      area #area_three {
        width: '5%'
        display: block
      }
      area #area_four {
        width: '14%'
        display: block
      }
      area #area_five_space {
        width: '11%'
        display: block
      }
      area #area_five {
        width: '5%'
        display: block
      }
      area #area_six {
        width: '16%'
        display: block
      }
    }
    tile text #textTile_01 {
      areaId: area_two
      value: "Response Rate"
      style {
        fontSize: 24
      }

    }

    tile value #valueTile_1 {
      areaId: area_two
      value: 100 * @cp.WFComplete / COUNT(:responseid)
      valueFormatter: percentNoDecimal
      style {
        fontSize: 40
        //fontWeight: bold
        color: #000000
        A {
        }

      }
      valueColorFormatter: dropOffDefaultFormatter
    }
    tile chartPlus #icon1 {
      areaId: area_one
      palette: icon_pie_palette
      style {
        height: 100px
      }
      chart pie {
        innerRadius: 30
        outerRadius: 45
        legendType: circle
      }
      series {
        label: "Responses"
        value: COUNT(:responseid) / count(:, true, "__top") * 100
        base: COUNT(:responseid)
        valueFormatter: statisticPercentsDefaultFormatter
      }
      category cut {
        value: :status
      }
      removeEmptyCategories: true


    }
    tile text #textTile_02 {
      areaId: area_four
      value: "Number Invited"
      style {
        fontSize: 24
        color: #000000
      }
    }
    tile value #valueTile_4 {
      areaId: area_four
      value: COUNT(:responseid)
      valueFormatter: bigNumberFormatter
      style {
        fontSize: 40
        color: #000000
      }
    }
    tile text #textTile_03 {
      areaId: area_six
      value: "Completed Surveys"
      style {
        fontSize: 24
      }
    }
    tile value #valueTile_3 {
      areaId: area_six
      value: @cp.WFComplete
      valueFormatter: bigNumberFormatter
      style {
        fontSize: 40
        color: #000000

      }
    }
    tile image #imageTile {
      areaId: area_three
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/file%20library%20test/RR_Invite.jpg"
    }
    tile image #imageTile_2 {
      areaId: area_five
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/file%20library%20test/RR_Complete.jpg"
    }
  }
  widget headline #summaryMTVPrimaryDimDonut {
    label: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.label
    description: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.description
    hide: @rollupMode.selected.mode != "rollup"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.infoText
          label: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {
        action navigate {
          navigateTo: orgDetails
        }
      }
    }

    cell: @dtEngagementSummary.m.data.main
    //CNJ126 replaced container
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      area #labelFirst {
        width: '29%'
        display: block
        paddingLeft: 15px
      }
      area #labelSecond {
        display: block
        width: '60%'
        paddingLeft: 60px
      }
      // area #labelThird {
      //   display: block
      //   width: '35%'
      //   paddingLeft: 30px
      // }
      area #left {
        width: '30%'
        height: 300px
        paddingLeft: 50px

        position: relative
        area #donut {
          position: absolute
        }
        area #center {
          position: absolute
        }
      }
      // area #legend {
      //   width: '15%'
      //   display: flex
      //   flexDirection: column
      //   alignItems: baseline
      // }


      area #right {
        width: '70%'
        display: block
        paddingLeft: 30px
        paddingBottom: 30px
      }
      area #legend {
        width: '100%'
        paddingLeft: 20px
        paddingBottom: 30px

      }
    }


    filter expression {
      value: .dimensions:id = "engagement"
    }
    tile text #textTile_3 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelFirst
      value: "Engagement Mean Score and Level Distribution"
    }
    tile text #textTile_4 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelSecond
      value: "Items Included in Your Engagement Score"

    }
    // tile text #textTile_5 {
    //   style {
    //     fontSize: 16px
    //     fontWeight: bold
    //   }
    //   areaId: labelThird
    //   value: "Items Included in Your Engagement Score"
    // }

    tile microchart #microchartTile_2 {
      areaId: donut
      value: @dtEngagementSummary.m.data.microchart.value
      microchart pie {
        donutWidth: 30%
        percentFormat: percentNoDecimal
        //CNJ126 legend
        legendType: diamond
        palette: engaged
      }
      style {
        width: "350px"
        height: "250px"
      }
      legend: bottomCenter

    }


    tile custom #customTile_2 {
      areaId: center
      expression #score {
        value: @cell.current
        valueFormatter: scoreFormatter
      }
      expression #change {
        value: @cell.change
        valueFormatter: scoreFormatter
      }
      expression #percentile {
        value: @dtEngagementSummary.m.data.benchmark.rank
        formatter: rankFormatter
      }
      expression #asteric {
        value: @cell.asteric//IIF(@cell.sig != 0, "*", " ")
      }
      expression #arrow {
        value: @cell.arrow//IIF(@cell.change > 0, "↑", IIF(change[] < 0, "↓", "-"))
      }
      expression #sigInfo {
        value: @cell.sigInfo// IIF(@cell.sig != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      formula #color {
        value: IIF(change[] > 0, IIF(@cell.sig != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(@cell.sig != 0, "#d02625", "Black"), "Black"))
      }
      formula #historyMean {
        value: @cell.current - @cell.change
        formatter: floatDefaultFormatter
      }
      //CNJ126 arrows edited formatstring
      formatString: '{score} <span style="color:{color}">{arrow}</span> {asteric}<span style="font-size: 16px; color:grey; display:block">{percentile} percentile</span>'
      tooltipFormatString: "<span style='font-size:40px'>{historyMean}</span><br>Mean Score for " + @surveyToCompareWith.selectedLabel + "<br><br><span style='font-size:30px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigInfo}"

      style {
        fontSize: 40px
        display: block
        textAlign: center
      }
    }

    //CNJ126 Tile legend  For different legends; try ● ■
     //but then you should also change legendtype on Key drivers, datagrids and tooltips
    tile custom #legend_1 {
      areaId: legend
      formatString: '<span style="color:#027580"> ✦ </span> Highly Engaged'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_2 {
      areaId: legend
      formatString: '<span style="color:#1BA583">✦ </span> Engaged'
      style {
        fontSize: 14
      }
    }
    tile custom #legend_3 {
      areaId: legend
      formatString: '<span style="color:#E69F0D">✦ </span> Neutral'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_4 {
      areaId: legend
      formatString: '<span style="color:#D02624">✦ </span> Disengaged'
      style {
        fontSize: 14
      }
    }

    // tile chartPlus #summaryMTVTrend {
    //   label: @widgetConfig.lookup.data.summaryMTVTrend.label
    //   description: @widgetConfig.lookup.data.summaryMTVTrend.description
    //   hide: @rollupMode.selected.mode != "rollup"
    //   areaId: middle

    //   scope filter {
    //     name: period
    //     value: AllPeriods
    //   }


    //   filter expression {
    //     value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    //   }
    //   category cut #periods {
    //     value: .reportHistory:trendYear
    //     sortBy: .reportHistory:trendYear
    //     sortOrder: ascending
    //   }

    //   series {
    //     label: ""
    //     value: parseInt("a")
    //     chart bar {
    //       legendType: none
    //     }
    //   }

    //   axis category {
    //     interval: preserveStartEnd
    //   }

    //   series #user {
    //     label: @rollupMode.selectedLabel
    //     value: :dimensionScore()
    //     chart line {
    //     }
    //   }
    //   series #entire {
    //     label: "Entire organization"
    //     scope reportingHierarchy {
    //       reportingHierarchy: unitHierarchy
    //       nodes: AllData
    //     }
    //     filter expression {
    //       value: _isNotNull(@unitHierarchy.source)
    //     }
    //     value: :dimensionScore()
    //     chart line {
    //     }
    //   }
    //   series #benchm {

    //     label: @defaultBenchmmark.selected.definitionName
    //     value: lookup value {
    //       source: benchmarks
    //       mapping value {
    //         value: @externalConfig.primaryDimensionId
    //         selector: bmValueCode
    //       }
    //       mapping value {
    //         value: @defaultBenchmmark.selected.definitionId
    //         selector: benchmarkDefinitionID
    //       }
    //       mapping header {
    //         header: periods
    //       //value: .reportHistory:trendYear
    //         selector: TrendYear
    //       }
    //       value: mean
    //       formatter: scoreFormatter
    //     }
    //     chart line {
    //     }
    //   }
    //   legend: rightMiddle
    //   axis primary {
    //   }

    //   axis secondary #secondaryAxis {
    //     hide: true
    //   }
    // }


    tile grid #gridTile_2 {

      areaId: right
      style {
        width: "100%"
      }
      showBullets: false

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }
      row #headerLabels {
        label: " "
        cell custom {
          row: headerLabels
          column: main
          formula #value {
            value: "Mean Score"
          }
          formatString: "<b>{value}</b>"
        }
      }
      cell custom { //Errors out if you put too many cells 
        row: headerLabels
        column: benchmark
        formula #value {
          value: "Percentile Rank"
        }
        formatString: "<b>{value}</b>"
      }
      row list #items {
        table: .items:
        value: answerText(.items:Id) //toText(.items:SequenceId) + ". " +
      }

      column cut #history {
        hide: true
        //categories: "'_1'"
        scope filter {
          name: period
          value: currentAndPrevious
        }
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :itemScore()
          }
          statistic mean #sig {
            testingType: T
            argument: numeric(.item_score:questionScoreValue)
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diffSum}"
          tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

        }
      }
      column #main {
        label: "Mean Score"
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #asteric {
            value: IIF(sig[column = /history.current] != 0, "*", " ")
          }
          formula #sigText {
            value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.1] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
          }
          formula #historyMean {
            value: score[column = /history.current] - diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }

          formatString: "<pre>{current}<span style='font-size:20px; color:{color};'>{arrow}</span>{asteric}</pre>"
          tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        }
      }
      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: :itemScore()
            formatter: rankFormatter
          }
          lookup value #mean {
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: mean
            formatter: scoreFormatter
          }
          formula #tooltip {
            value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>Benchmark Mean Value: " + mean[], "too few responses")
            //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
          }
          formatString: "{rank}"
          tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
    //          tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

        }
      }
    }
    size: halfwidth
  }

  widget chart #summaryMTVTrend {
    label: @widgetConfig.lookup.data.summaryMTVTrend.label
    description: @widgetConfig.lookup.data.summaryMTVTrend.description
    hide: @rollupMode.selected.mode != "rollup"
    //animation: true
  // chart line #barChart {
  //   lineType: monotone
  //   lineWidth: 2
  //   dotSize: 5
  // }

    series {
      label: " "
      value: parseInt("a")
      chart bar {
        legendType: none
      }
    }
    series #user {
      label: @rollupMode.selectedLabel
      value: :dimensionScore()
      chart line {
        lineType: monotone
      }
    }


    scope filter {
      name: period
      value: AllPeriods
    }

    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }
    category cut #periods {
      value: .reportHistory:trendYear
      sortBy: .reportHistory:trendYear
      sortOrder: ascending
    }
    axis category {
      interval: preserveStartEnd
    }

    series #entire {
      label: "Overall Organization"
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      value: :dimensionScore()
      chart line {
        lineType: monotone
      }
    }

    series #benchmark {
      label: @defaultBenchmmark.selected.definitionName
      value: lookup value {
        source: benchmarks
        mapping value {
          value: @externalConfig.primaryDimensionId
          selector: bmValueCode
        }
        mapping value {
          value: @defaultBenchmmark.selected.definitionId
          selector: benchmarkDefinitionID
        }
        mapping header {
          header: periods
          selector: TrendYear
        }
        value: mean
        formatter: scoreFormatter
      }
      chart line {
        lineType: monotone
      }
      legend: rightMiddle
      axis primary {
      }
      axis secondary #secondaryAxis {
        hide: true
      }
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: medium
  } //here   
  widget headline #summaryMTVLargeGroups_Eng {

    size: large
    label: @widgetConfig.lookup.data.summaryMTVLargeGroups_Eng.label
    description: @widgetConfig.lookup.data.summaryMTVLargeGroups_Eng.description
    hide: @rollupMode.selected.mode != "rollup"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected
      label: "The number of responses for your team is below the minimum theshold required to display results."
    }
    toolbar {
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVLargeGroups_Eng.infoText
          label: @widgetConfig.lookup.data.summaryMTVLargeGroups_Eng.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }
      button #navigate {
        action navigate {
          navigateTo: page_5
        }
          // action setSelector {
          //   value: Engagement
          //    select: @dimensionsSelector2
          // }
      }
    }

    //CNJ126 padding botttom
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      area #donuts {
        width: '100%'
        display: flex
        paddingLeft: 30px
        paddingBottom: 30px
        justifyContent: "center"//"space-evenly"
      }
      area #legend {
        width: '100%'
        paddingLeft: 20px
        paddingBottom: 30px

      }
    }


    tile set #setTile_2 {
      areaId: donuts

      //CNJ126 tileset switch container flex with grid
      container: container grid {
        rows: 'A A A A A'
        justifyContent: spaceEvenly

      }
      /* container: container flex {
        flexDirection: row
        flexWrap: wrap
      } */
      itemContainer: container flex {
        flexDirection: column
          // backgroundColor: yellow
        width: 300px
          //display: flex

        area #label {
          height: 50px
          display: block
        }
        area #respondents {
            // height: 10px
          display: block
        }
        area #main {
          //  width: 500px
          //  height: 500px
            // backgroundColor: orange
          position: relative
          area #donut {
              // backgroundColor: green
              //position: absolute
              // top: "50%"
              // left: "50%"
              // transform: "translate(-50%, -50%)"
          }
          area #center {
              // backgroundColor: orange
            position: absolute
              // top: "50%"
              // left: "50%"
              // transform: "translate(-50%, -50%)"
          }
        }
      }

      breakdownBy inlineData {
        value: @dtEngagementNodes.m.data
      }

      tile text {
        areaId: label
        value: this.nodeLabel.value
        style {
          fontSize: 15px
          //fontWeight: bold
        }
      }
      tile value {
        areaId: respondents
        value: this.base.value
        formatString: "{value} Responses"
        style {
          fontSize: 16px
        }
      }

      tile microchart {
        areaId: donut
        value: this.microchart.value
        microchart pie {
          donutWidth: 30px
          palette: engaged
          valuePosition: outer
          percentFormat: percentNoDecimal

        }
        style {
          height: 205px
          width: 260px
            // paddingBottom:25px

        }
      }


      tile custom #customTile_2 {
        areaId: center
        expression #score {
          value: this.main.score
          valueFormatter: scoreFormatter
        }
        expression #change {
          value: this.main.change
          valueFormatter: scoreFormatter
        }
        expression #percentile {
          value: this.benchmark.rank
          formatter: rankFormatter
        }
        expression #asteric {
          value: this.main.asteric//IIF(this.main.sig != 0, "*", " ")
        }
        expression #arrow {
          value: this.main.arrow//IIF(this.main.change > 0, "↑", IIF(this.main.change < 0, "↓", "-"))
        }
        expression #sigInfo {
          value: this.main.sigInfo//IIF(this.main.sig != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        expression #label {
          value: this.main.label
        }
        expression #color {
          value: this.main.color
        }
        expression #historyMean {
          value: this.main.historyMean
        }
      //CNJ126 arrows edited formatstring
        formatString: '<span style="font-size: 30px; display:block">{score} <span style="color:{color}">{arrow}</span> {asteric}</span><span style="font-size: 14px; color:grey; display:block">{percentile} Percentile</span>'
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigInfo}"


          // formatString: '{score} {arrow} {asteric}<span style="font-size: 20px; display:block">{percentile} percentile</span>'
          // tooltipFormatString: "change {change} vs {}label}" + "<br/>{sigInfo}"

        style {
          fontSize: 40px
          display: block
          textAlign: center
        }
      }



    }

    tile custom #legend_1 {
      areaId: legend
      formatString: '<span style="color:#027580"> ✦ </span> Highly Engaged'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_2 {
      areaId: legend
      formatString: '<span style="color:#1BA583">✦ </span> Engaged'
      style {
        fontSize: 14
      }
    }
    tile custom #legend_3 {
      areaId: legend
      formatString: '<span style="color:#E69F0D">✦ </span> Neutral'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_4 {
      areaId: legend
      formatString: '<span style="color:#D02624">✦ </span> Disengaged'
      style {
        fontSize: 14
      }
    }

  }

  // widget headline #summaryMTVLeaderIndex {
  //   label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
  //   description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
  //   hide: @rollupMode.selected.mode != "rollup"

  //   suppressRule {
  //     criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected //when
  //     label: "The number of responses for your team is below the minimum threshold." //what to display
  //   }
  //   toolbar { // This 
  //     button #infobox {
  //       action showInfobox {
  //         size: large
  //         info: @widgetConfig.lookup.data.summaryMTVLeaderIndex.infoText
  //         label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
  //       }
  //     }
  //     button #export {
  //       action export {
  //         format: png
  //       }
  //     }

  //     button #navigate {

  //       action navigate {
  //         navigateTo: orgDetails
  //       }

  //     }
  //   }


  //   // suppressRule {
  //   //   criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected
  //   //   label: "The number of responses for your team is below the minimum threshold required to display results."
  //   // }

  //   cell: @dtEngagementSummary.m.data.main
  //   container: container flex {
  //     flexDirection: row
  //     flexWrap: wrap
  //     //Area for labels
  //     area #labelFirst {
  //       width: '29%'
  //       display: block
  //       paddingLeft: 40px
  //       // paddingBottom:20px
  //     }
  //     area #labelSecond {
  //       width: '30%'
  //       display: block
  //       paddingLeft: 30px
  //     }
  //     area #labelThird {
  //       display: block
  //       width: '40%'

  //     }
  //     // area #labelFourth {
  //     //   display: block
  //     //   width: '7%'
  //     //   // paddingLeft: 34px
  //     // }
  //     //Area for charts and tables
  //     area #left {
  //       width: "25%"
  //     }
  //     area #middle {
  //       width: "30%"
  //       paddingLeft: 40px
  //       height: 400px
  //       position: relative
  //       area #donut {
  //         position: absolute
  //       }
  //       area #center {
  //         position: absolute
  //       }
  //     }
  //     area #right {
  //       width: "40%"
  //       //paddingLeft: 40px
  //     }
  //   }


  //   filter expression {
  //     value: .dimensions:id = "leaderindex"
  //   }

  //   //Text Tiles for Headers
  //   tile text #textTile_2 {
  //     style {
  //       fontSize: 16px
  //       fontWeight: bold
  //     }
  //     areaId: labelFirst
  //     value: "Overall Leader Index for Your Team"
  //   }
  //   tile text #textTile_3 {
  //     style {
  //       fontSize: 16px
  //       fontWeight: bold
  //     }
  //     areaId: labelSecond
  //     value: "Group Distribution by Leader Index Score"
  //   }
  //   tile text #textTile_4 {
  //     style {
  //       fontSize: 16px
  //       fontWeight: bold
  //     }
  //     areaId: labelThird
  //     value: "Items Included in Your Leader Index"
  //   }
  //   // tile text #textTile_5 {
  //   //   style {
  //   //     fontSize: 18px
  //   //     fontWeight: bold
  //   //   }
  //   //   areaId: labelThird
  //   //   value: "Mean Score"
  //   // }
  //   // tile text #textTile_6 {
  //   //   style {
  //   //     fontSize: 18px
  //   //     fontWeight: bold
  //   //   }
  //   //   areaId: labelFourth
  //   //   value: "Percentile Rank"
  //   // }

  //   //Chart and Table Tiles
  //   tile custom #leaderindex {
  //     expression #score {
  //       value: :dimensionScore()
  //       valueFormatter: scoreFormatter
  //     }
  //     expression #color {
  //       value: IIF(:dimensionScore() >= 4, "#1FA583", IIF(:dimensionScore() <= 2.5, "#D02525", "#E79F0B"))
  //     }
  //     expression #label {
  //       value: IIF(:dimensionScore() >= 4, "High", IIF(:dimensionScore() <= 2.5, "#D02525", "Moderate"))

  //     }
  //     expression #description {
  //       value: IIF(:dimensionScore() >= 4, "Group is ready to have improvement planning discussions with their direct leader.", IIF(:dimensionScore() <= 2.5, "Focus should be placed on building relationships between direct leader and team prior to improvement planning.", "Group may be ready for improvement planning discussions, but the direct leader may benefit from additional guidance."))
  //     }
  //   //cb here
  //     areaId: left

  //     formatString: '<span style= "margin-left:200px;"><span style="font-size:60px";> {score}</span><br><span style="font-size:40px; margin-left:210px; color:{color};">{label}</span><br><br><p style="font-size:16px; margin-left:30px;">{description}</p>'

  //   }
  //   tile chartPlus #t1 {
  //     // filter expression {
  //     //   value: :combined_sourceid = "p494984785246"
  //     // }
  //     areaId: donut
  //     style {
  //       width: 350px
  //       paddingBottom: 10px
  //     }
  //     //test if palette work
  //     // palette: posNeuNeg

  //     axis primary #primaryAxis {
  //       hide: true
  //     }
  //     chartMargin {
  //       top: 40
  //     }
  //     series {
  //       label: "Responses"
  //       //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
  //       value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
  //       // removeEmptySeries: true
  //       base: count(unitHierarchy:)
  //       chart bar {
  //         // mode: stacked
  //         showBase: true
  //         valueLabel: "Groups"
  //         valuePosition: outer
  //       }
  //       format: percentNoDecimal
  //     }
  //     category cut {
  //       //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
  //       value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
  //       palette: LIpalette

  //     }
  //   }




  //   tile grid #gridTile_2 {

  //     areaId: right
  //     style {
  //       width: "100%"
  //     }
  //     showBullets: false

  //     suppression recordsBase {
  //       threshold: @suppressionThreshold.selected
  //     }

  //     row #headerLabels {
  //       label: " "
  //       cell custom {
  //         row: headerLabels
  //         column: main
  //         formula #value {
  //           value: "Mean Score"
  //         }
  //         formatString: "<b>{value}</b>"
  //       }
  //     }
  //     cell custom { //Errors out if you put too many cells 
  //       row: headerLabels
  //       column: benchmark
  //       formula #value {
  //         value: "Percentile Rank"
  //       }
  //       formatString: "<b>{value}</b>"
  //     }
  //     row list #items {
  //       table: .items:
  //       value: answerText(.items:Id) //toText(.items:SequenceId) + ". " + 
  //     }

  //     column cut #history {
  //       hide: true
  //       //categories: "'_1'"
  //       scope filter {
  //         name: period
  //         value: currentAndPrevious
  //       }
  //       total: none
  //       value: .reportHistory:historyTypeCode
  //       cell custom {
  //         expression #score {
  //           value: :itemScore()
  //         }
  //         statistic mean #sig {
  //           testingType: T
  //           argument: numeric(.item_score:questionScoreValue)
  //           compare: next
  //         }
  //         formula #diff {
  //           value: score[column = %.current] - score[]
  //         }
  //         formula #diffSum {
  //           value: sum(diff[column = %.*])
  //         }
  //         formatString: "{score} [{sig}] {diffSum}"
  //         tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
  //       }
  //     }
  //     column #main {
  //       cell custom {
  //         formula #current {
  //           value: score[column = /history.current]
  //         }
  //         formula #change {
  //           value: diffSum[column = /history.current]
  //           formatter: floatDefaultFormatter
  //         }
  //         formula #arrow {
  //           //CNJ126 arrows ↑↓ or  ↑ ↓
  //           value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
  //         }
  //         formula #asteric {
  //           value: IIF(sig[column = /history.current] != 0, "*", " ")
  //         }
  //         formula #sigText {
  //           value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
  //         }
  //         formula #color {
  //           value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
  //         }
  //         formula #historyMean {
  //           value: score[column = /history.current] - diffSum[column = /history.current]
  //           formatter: floatDefaultFormatter
  //         }
  //         formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
  //         tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

  //       }
  //     }
  //     column #benchmark {
  //       cell custom {
  //         lookup rank #rank {
  //           takeInArray: Per
  //           mode percentile {
  //           }
  //           source: benchmarks
  //           mapping header {
  //             header: items
  //             selector: bmValueCode
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.definitionId
  //             selector: BenchmarkDefinitionId
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.periodId
  //             selector: TrendYear
  //           }
  //           value: :itemScore()
  //           formatter: rankFormatter
  //         }
  //         lookup value #mean {
  //           source: benchmarks
  //           mapping header {
  //             header: items
  //             selector: bmValueCode
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.definitionId
  //             selector: BenchmarkDefinitionId
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.periodId
  //             selector: TrendYear
  //           }
  //           value: mean
  //           formatter: scoreFormatter
  //         }
  //         formula #tooltip {
  //           value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
  //           //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
  //         }
  //         formatString: "{rank}"
  //         tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
  //   //tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

  //       }
  //     }
  //   }
  //   size: large
  // }

  widget headline #summaryMTVLeaderIndex {
    label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
    description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
    hide: @rollupMode.selected.mode != "rollup"

    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold." //what to display
    }
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVLeaderIndex.infoText
          label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: orgDetails
        }

      }
    }


    // suppressRule {
    //   criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected
    //   label: "The number of responses for your team is below the minimum threshold required to display results."
    // }

    cell: @dtEngagementSummary.m.data.main
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      //Area for labels
      area #labelFirst {
        width: '40%'
        display: block
        paddingLeft: 15px
      }
      // area #labelSecond {
      //   width: '30%'
      //   display: block
      //   //paddingLeft: 30px
      // }
      area #labelThird {
        display: block
        width: '50%'
        // paddingLeft: 10px
      }

      area #left {
        width: '35%'
        //display: block
        // height:300px
      }
      // area #middle {
      //   width: '30%'
      //   paddingLeft: 15px
      //   display: block
      //   height: 300px
      //   /* position: relative
      //   area #donut {
      //     position: absolute
      //   } */
      //   /* area #center {
      //     position: absolute
      //   } */
      // }
      area #right {
        width: '60%'
        display: block

      }
    }


    filter expression {
      value: .dimensions:id = "leaderindex"
    }

    //Text Tiles for Headers
    tile text #textTile_2 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelFirst
      value: "Overall Leader Index for Your Team"
    }
    // tile text #textTile_3 {
    //   style {
    //     fontSize: 16px
    //     fontWeight: bold
    //   }
    //   areaId: labelSecond
    //   value: "Group Distribution by Leader Index Score"
    // }
    tile text #textTile_4 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelThird
      value: "Items Included in Your Leader Index"
    }
    // tile text #textTile_5 {
    //   style {
    //     fontSize: 18px
    //     fontWeight: bold
    //   }
    //   areaId: labelThird
    //   value: "Mean Score"
    // }
    // tile text #textTile_6 {
    //   style {
    //     fontSize: 18px
    //     fontWeight: bold
    //   }
    //   areaId: labelFourth
    //   value: "Percentile Rank"
    // }

    //Chart and Table Tiles
    tile custom #leaderindex {

      areaId: left
      expression #score {
        value: @cell.current
        valueFormatter: scoreFormatter
      }
      expression #change {
        value: @cell.change
        valueFormatter: scoreFormatter
      }
      expression #percentile {
        value: @dtEngagementSummary.m.data.benchmark.rank
        formatter: rankFormatter
      }
      expression #asteric {
        value: @cell.asteric//IIF(@cell.sig != 0, "*", " ")
      }
      expression #arrow {
        value: @cell.arrow//IIF(@cell.change > 0, "↑", IIF(change[] < 0, "↓", "-"))
      }
      expression #sigInfo {
        value: @cell.sigInfo// IIF(@cell.sig != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      formula #arrowColor {
        value: IIF(change[] > 0, IIF(@cell.sig != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(@cell.sig != 0, "#d02625", "Black"), "Black"))
      }
      formula #historyMean {
        value: @cell.current - @cell.change
        formatter: floatDefaultFormatter
      }
      // expression #score {
      //   value: :dimensionScore()
      //   valueFormatter: scoreFormatter
      // }
      expression #color {
        value: IIF(@cell.current >= 4, "#1FA583", IIF(@cell.current <= 2.5, "#D02525", "#E79F0B"))
      }
      expression #label {
        value: IIF(@cell.current >= 4, "High", IIF(@cell.current <= 2.5, "#D02525", "Moderate"))

      }
      //     formula #current {
      //       value: score[column = /history.current]
      //     }
      //     formula #change {
      //       value: diffSum[column = /history.current]
      //       formatter: floatDefaultFormatter
      //     }
      //     formula #arrow {
      //       //CNJ126 arrows ↑↓ or  ↑ ↓
      //       value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
      //     }
      //     formula #asteric {
      //       value: IIF(sig[column = /history.current] != 0, "*", " ")
      //     }
      formula #sigText {
        value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      //               formula #arrowColor {
      //       value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
      //     }
      //     formula #historyMean {
      //       value: score[column = /history.current] - diffSum[column = /history.current]
      //       formatter: floatDefaultFormatter
      //     }

      expression #description {
        value: IIF(:dimensionScore() >= 4, "Group is ready to have improvement planning discussions with their direct leader.", IIF(:dimensionScore() <= 2.5, "Focus should be placed on building relationships between direct leader and team prior to improvement planning.", "Group may be ready for improvement planning discussions, but the direct leader may benefit from additional guidance."))
      }
      //cb here

      formatString: '<span style= "margin-left:80px;font-size:60px"> {score}</span><span style ="color:{arrowColor}">{arrow}</span><br><span style="font-size:40px; margin-left:95px; color:{color};">{label}</span><br><br><p style="font-size:16px; margin-left:10px;">{description}</p>'
      tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {arrowColor};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

    }
    // tile chartPlus #t1 {
    //   // filter expression {
    //   //   value: :combined_sourceid = "p494984785246"
    //   // }
    //   areaId: middle
    //   style {
    //     width: 500px
    //     height: 260px
    //     //paddingBottom: 10px
    //   }
    //   //test if palette work
    //   // palette: posNeuNeg

    //   axis primary #primaryAxis {
    //     hide: true
    //   }
    //   chartMargin {
    //     top: 40
    //   }
    //   series {
    //     label: "Responses"
    //     //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
    //     value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
    //     // removeEmptySeries: true
    //     base: count(unitHierarchy:)
    //     chart bar {
    //       // mode: stacked
    //       showBase: true
    //       valueLabel: "Groups"
    //       valuePosition: outer
    //     }
    //     format: percentNoDecimal
    //   }
    //   category cut {
    //     //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
    //     value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
    //     palette: LIpalette

    //   }
    // }




    tile grid #gridTile_2 {

      areaId: right
      style {
        width: "100%"
      }
      showBullets: false

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }

      row #headerLabels {
        label: " "
        cell custom {
          row: headerLabels
          column: main
          formula #value {
            value: "Mean Score"
          }
          formatString: "<b>{value}</b>"
        }
      }
      cell custom { //Errors out if you put too many cells 
        row: headerLabels
        column: benchmark
        formula #value {
          value: "Percentile Rank"
        }
        formatString: "<b>{value}</b>"
      }
      row list #items {
        table: .items:
        value: answerText(.items:Id) //toText(.items:SequenceId) + ". " + 
      }

      column cut #history {
        hide: true
        //categories: "'_1'"
        scope filter {
          name: period
          value: currentAndPrevious
        }
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :itemScore()
          }
          statistic mean #sig {
            testingType: T
            argument: numeric(.item_score:questionScoreValue)
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diffSum}"
          tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
        }
      }
      column #main {
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #asteric {
            value: IIF(sig[column = /history.current] != 0, "*", " ")
          }
          formula #sigText {
            value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
          }
          formula #historyMean {
            value: score[column = /history.current] - diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }

          formatString: "<pre>{current}<span style='color:{color};font-size:20px;'>{arrow}</span>{asteric}</pre>"
          tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        }
      }
      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: :itemScore()
            formatter: rankFormatter
          }
          lookup value #mean {
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: mean
            formatter: scoreFormatter
          }
          formula #tooltip {
            value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
            //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
          }
          formatString: "{rank}"
          tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
    //tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

        }
      }
    }
    size: medium
  }

  widget chart #summaryMTVLeaderIndexChart {
    label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
    description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
    hide: @rollupMode.selected.mode != "rollup"
    st {
    }
    series {
      label: "Responses"
        //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
      value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
        // removeEmptySeries: true
      base: count(unitHierarchy:)
      chart bar {
          // mode: stacked
        showBase: true
        valueLabel: "Groups"
        valuePosition: outer
        maxBarSize: 125

      }
      format: percentNoDecimal
    }
    category cut {
        //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
      value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
      palette: LIpalette

    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {

      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: medium
  }


  widget dataGrid #summaryMTVKeyDrivers {
    label: @widgetConfig.lookup.data.summaryMTVKeyDrivers.label
    description: @widgetConfig.lookup.data.summaryMTVKeyDrivers.description
    size: medium
    hide: @rollupMode.selected.mode != "rollup"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVKeyDrivers.infoText
          label: @widgetConfig.lookup.data.summaryMTVKeyDrivers.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/score100"
      sortOrder: descending
      takeTop: 6
    }


   //filterexpression{ value: .dimension_score:dg1_dimensionScore = "Standard_3" }			

    row cut #itemsRow {
      total: none
      value: .item_score:dg1_questionScore
      filter expression {
        value: .scaled_items:includeKD
      }

    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:)
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint

        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }
    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }
    }

    column #gpr {
      label: "Percentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }



  widget dataGrid #summaryMTVTopPerform {
    label: @widgetConfig.lookup.data.summaryMTVTopPerform.label
    description: @widgetConfig.lookup.data.summaryMTVTopPerform.description
    size: medium
    hide: @rollupMode.selected.mode != "rollup"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVTopPerform.infoText
          label: @widgetConfig.lookup.data.summaryMTVTopPerform.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/gpr"
      sortOrder: descending
      takeTop: 5
    }

    row cut #itemsRow {
      total: none
      value: .item_score:dg1_questionScore


    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:)
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint
        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }

    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }


    }



    column #gpr {
      label: "Precentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }
  widget chart #keyDemoChartTop {
    label: "Top Performing Demographic Groups"// @widgetConfig.lookup.data.summaryMTVKeyDemo.label
    description: @widgetConfig.lookup.data.summaryMTVKeyDemo.description
    size: medium
    layout: vertical
    legend: bottomCenter
    hide: @rollupMode.selected.mode != "rollup"
    axis category {
      textSize: 150

    }


    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }

    category cutByMulti {
      value: :keyDemoCalc
      sortBy: "/score"
      sortOrder: descending
      takeTop: 3
      //total: none

    }
    // series {
    //   label: @defaultBenchmmark.selectedLabel
    //   value: lookup value {
    //     source: benchmarks
    //     mapping value {
    //       value: @externalConfig.primaryDimensionId
    //       selector: bmValueCode
    //     }
    //     mapping value {
    //       value: @defaultBenchmmark.selected.definitionId
    //       selector: BenchmarkDefinitionId
    //     }
    //     mapping value {
    //       value: @defaultBenchmmark.selected.periodId
    //       selector: TrendYear
    //     }
    //     value: mean
    //     formatter: scoreFormatter
    //   }

    // }

    series #score {
      label: "Engagement mean score"
      value: IIF(count(:) > 5 AND count(:) / count(:, true, "__top") > 0.03, :dimensionScore())

    }

    axis primary #primaryAxis {
      maxValue: 5
      minValue: 0
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    significanceTesting: true
  }

  widget chart #keyDemoChartBottom {
    label: "Bottom Performing Demographic Groups"//@widgetConfig.lookup.data.summaryMTVKeyDemo.label
    description: @widgetConfig.lookup.data.summaryMTVKeyDemo.description
    size: medium
    layout: vertical
    legend: bottomCenter
    hide: @rollupMode.selected.mode != "rollup"
    axis category {
      textSize: 150
    }

    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }

    category cutByMulti {
      value: :keyDemoCalc
      sortBy: "/score"
      sortOrder: ascending
      takeTop: 3
      //total: none

    }
    // series {
    //   label: @defaultBenchmmark.selectedLabel
    //   value: lookup value {
    //     source: benchmarks
    //     mapping value {
    //       value: @externalConfig.primaryDimensionId
    //       selector: bmValueCode
    //     }
    //     mapping value {
    //       value: @defaultBenchmmark.selected.definitionId
    //       selector: BenchmarkDefinitionId
    //     }
    //     mapping value {
    //       value: @defaultBenchmmark.selected.periodId
    //       selector: TrendYear
    //     }
    //     value: mean
    //     formatter: scoreFormatter
    //   }

    // }

    series #score {
      label: "Engagement mean score"
      value: IIF(count(:) > 5 AND count(:) / count(:, true, "__top") > 0.03, :dimensionScore())


    }

    axis primary #primaryAxis {
      maxValue: 5
      minValue: 0
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    removeEmptyCategories: true
  }


  widget dataGrid #summaryMTVAddDimensions {
    label: @widgetConfig.lookup.data.summaryMTVAddDimensions.label
    description: @widgetConfig.lookup.data.summaryMTVAddDimensions.description
    hide: @rollupMode.selected.mode != "rollup"
    size: large
    filter expression {
      value: .dimensions:includeHXWidget
    }
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVAddDimensions.infoText
          label: @widgetConfig.lookup.data.summaryMTVAddDimensions.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }

    row list #dimensions {
      table: .dimensions:
      value: .dimensions:id
      total: none
    }

    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :dimensionScore()
        }
        statistic mean #sig {
          testingType: T
          argument: .dimension_score:dimensionScoreValue
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
      }
    }
    // column #recoding {
    //   label: " "
    //   cell custom {
    //     expression #type {
    //       value: ToText(.dimensions:id)
    //     }
    //     formula #teamIndex {
    //         //later should be recoce()
    //       value: IIF(value[column = /history.current] >= @externalConfig.teamIndex1, "TI-1", IIF(score[column = /history.current] < @externalConfig.teamIndex2, "TI-3", "TI-2"))
    //     }
    //     formula #team {
    //       value: IIF(type[] = "teamindex", teamIndex[])
    //     }

    //     formatString: "{team}"
    //   }
    // }
    column #main {
      label: "Mean score"
      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          //CNJ126 arrows ↑↓ or  ↑ ↓
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='font-size: 20px; color:{color};'>{arrow}</span>{asteric}</pre>"//To add Astric: 
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        // tooltipFormatString: "<b style='font-size:20px'>{historyMean}</b><br>Historical Mean Score" + "<br><b style='font-size:20px'>{change}</b><br> vs " + @surveyToCompareWith.selectedLabel + "<br><span style='  height: 25px;  width: 25px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }
    column #benchmark {
      label: "Percentile"
      cell custom {
        lookup rank #rank {
          takeInArray: Per
          mode percentile {
          }
          source: benchmarks
          mapping header {
            header: dimensions
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :dimensionScore()
          formatter: rankFormatter
        }
        lookup value #mean {
          source: benchmarks
          mapping header {
            header: dimensions
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: mean
          formatter: scoreFormatter
        }
        formula #tooltip {
          value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
        }
        formatString: "{rank}"
        tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>" + @defaultBenchmmark.selectedLabel + " Mean Score "
      }
    }
    column #recoding {
      label: " "
      sortable: false
      cell custom {
        formatString: " "
      }
    }

  }

  widget headline #summaryDRPrimaryDim {
    label: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.label
    description: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.description
    hide: @rollupMode.selected.mode != "direct"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.infoText
          label: @widgetConfig.lookup.data.summaryMTVPrimaryDimDonut.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {
        action navigate {
          navigateTo: orgDetails
        }
      }
    }

    cell: @dtEngagementSummary.m.data.main
    //CNJ126 replaced container
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      area #labelFirst {
        width: '29%'
        display: block
        paddingLeft: 15px
      }
      area #labelSecond {
        display: block
        width: '60%'
        paddingLeft: 60px
      }
      // area #labelThird {
      //   display: block
      //   width: '35%'
      //   paddingLeft: 30px
      // }
      area #left {
        width: '30%'
        height: 300px
        paddingLeft: 50px

        position: relative
        area #donut {
          position: absolute
        }
        area #center {
          position: absolute
        }
      }
      // area #legend {
      //   width: '15%'
      //   display: flex
      //   flexDirection: column
      //   alignItems: baseline
      // }


      area #right {
        width: '70%'
        display: block
        paddingLeft: 30px
        paddingBottom: 30px
      }
      area #legend {
        width: '100%'
        paddingLeft: 20px
        paddingBottom: 30px

      }
    }


    filter expression {
      value: .dimensions:id = "engagement"
    }
    tile text #textTile_3 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelFirst
      value: "Engagement Mean Score and Level Distribution"
    }
    tile text #textTile_4 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelSecond
      value: "Items Included in Your Engagement Score"

    }
    // tile text #textTile_5 {
    //   style {
    //     fontSize: 16px
    //     fontWeight: bold
    //   }
    //   areaId: labelThird
    //   value: "Items Included in Your Engagement Score"
    // }

    tile microchart #microchartTile_2 {
      areaId: donut
      value: @dtEngagementSummary.m.data.microchart.value
      microchart pie {
        donutWidth: 30%
        percentFormat: percentNoDecimal
        //CNJ126 legend
        legendType: diamond
        palette: engaged
      }
      style {
        width: "350px"
        height: "250px"
      }
      legend: bottomCenter

    }


    tile custom #customTile_2 {
      areaId: center
      expression #score {
        value: @cell.current
        valueFormatter: scoreFormatter
      }
      expression #change {
        value: @cell.change
        valueFormatter: scoreFormatter
      }
      expression #percentile {
        value: @dtEngagementSummary.m.data.benchmark.rank
        formatter: rankFormatter
      }
      expression #asteric {
        value: @cell.asteric//IIF(@cell.sig != 0, "*", " ")
      }
      expression #arrow {
        value: @cell.arrow//IIF(@cell.change > 0, "↑", IIF(change[] < 0, "↓", "-"))
      }
      expression #sigInfo {
        value: @cell.sigInfo// IIF(@cell.sig != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      formula #color {
        value: IIF(change[] > 0, IIF(@cell.sig != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(@cell.sig != 0, "#d02625", "Black"), "Black"))
      }
      formula #historyMean {
        value: @cell.current - @cell.change
        formatter: floatDefaultFormatter
      }
      //CNJ126 arrows edited formatstring
      formatString: '{score} <span style="color:{color}">{arrow}</span> {asteric}<span style="font-size: 16px; color:grey; display:block">{percentile} percentile</span>'
      tooltipFormatString: "<span style='font-size:40px'>{historyMean}</span><br>Mean Score for " + @surveyToCompareWith.selectedLabel + "<br><br><span style='font-size:30px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigInfo}"

      style {
        fontSize: 40px
        display: block
        textAlign: center
      }
    }

    //CNJ126 Tile legend  For different legends; try ● ■
     //but then you should also change legendtype on Key drivers, datagrids and tooltips
    tile custom #legend_1 {
      areaId: legend
      formatString: '<span style="color:#027580"> ✦ </span> Highly Engaged'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_2 {
      areaId: legend
      formatString: '<span style="color:#1BA583">✦ </span> Engaged'
      style {
        fontSize: 14
      }
    }
    tile custom #legend_3 {
      areaId: legend
      formatString: '<span style="color:#E69F0D">✦ </span> Neutral'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_4 {
      areaId: legend
      formatString: '<span style="color:#D02624">✦ </span> Disengaged'
      style {
        fontSize: 14
      }
    }

    // tile chartPlus #summaryMTVTrend {
    //   label: @widgetConfig.lookup.data.summaryMTVTrend.label
    //   description: @widgetConfig.lookup.data.summaryMTVTrend.description
    //   hide: @rollupMode.selected.mode != "rollup"
    //   areaId: middle

    //   scope filter {
    //     name: period
    //     value: AllPeriods
    //   }


    //   filter expression {
    //     value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    //   }
    //   category cut #periods {
    //     value: .reportHistory:trendYear
    //     sortBy: .reportHistory:trendYear
    //     sortOrder: ascending
    //   }

    //   series {
    //     label: ""
    //     value: parseInt("a")
    //     chart bar {
    //       legendType: none
    //     }
    //   }

    //   axis category {
    //     interval: preserveStartEnd
    //   }

    //   series #user {
    //     label: @rollupMode.selectedLabel
    //     value: :dimensionScore()
    //     chart line {
    //     }
    //   }
    //   series #entire {
    //     label: "Entire organization"
    //     scope reportingHierarchy {
    //       reportingHierarchy: unitHierarchy
    //       nodes: AllData
    //     }
    //     filter expression {
    //       value: _isNotNull(@unitHierarchy.source)
    //     }
    //     value: :dimensionScore()
    //     chart line {
    //     }
    //   }
    //   series #benchm {

    //     label: @defaultBenchmmark.selected.definitionName
    //     value: lookup value {
    //       source: benchmarks
    //       mapping value {
    //         value: @externalConfig.primaryDimensionId
    //         selector: bmValueCode
    //       }
    //       mapping value {
    //         value: @defaultBenchmmark.selected.definitionId
    //         selector: benchmarkDefinitionID
    //       }
    //       mapping header {
    //         header: periods
    //       //value: .reportHistory:trendYear
    //         selector: TrendYear
    //       }
    //       value: mean
    //       formatter: scoreFormatter
    //     }
    //     chart line {
    //     }
    //   }
    //   legend: rightMiddle
    //   axis primary {
    //   }

    //   axis secondary #secondaryAxis {
    //     hide: true
    //   }
    // }


    tile grid #gridTile_2 {

      areaId: right
      style {
        width: "100%"
      }
      showBullets: false

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }
      row #headerLabels {
        label: " "
        cell custom {
          row: headerLabels
          column: main
          formula #value {
            value: "Mean Score"
          }
          formatString: "<b>{value}</b>"
        }
      }
      cell custom { //Errors out if you put too many cells 
        row: headerLabels
        column: benchmark
        formula #value {
          value: "Percentile Rank"
        }
        formatString: "<b>{value}</b>"
      }
      row list #items {
        table: .items:
        value: answerText(.items:Id) //toText(.items:SequenceId) + ". " +
      }

      column cut #history {
        hide: true
        //categories: "'_1'"
        scope filter {
          name: period
          value: currentAndPrevious
        }
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :itemScore()
          }
          statistic mean #sig {
            testingType: T
            argument: numeric(.item_score:questionScoreValue)
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diffSum}"
          tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

        }
      }
      column #main {
        label: "Mean Score"
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #asteric {
            value: IIF(sig[column = /history.current] != 0, "*", " ")
          }
          formula #sigText {
            value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.1] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
          }
          formula #historyMean {
            value: score[column = /history.current] - diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }

          formatString: "<pre>{current}<span style='font-size:20px; color:{color};'>{arrow}</span>{asteric}</pre>"
          tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        }
      }
      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: :itemScore()
            formatter: rankFormatter
          }
          lookup value #mean {
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: mean
            formatter: scoreFormatter
          }
          formula #tooltip {
            value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>Benchmark Mean Value: " + mean[], "too few responses")
            //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
          }
          formatString: "{rank}"
          tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
    //          tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

        }
      }
    }
    size: halfwidth
  }

  widget chart #summaryDRTrend {
    label: @widgetConfig.lookup.data.summaryDRTrend.label
    description: @widgetConfig.lookup.data.summaryDRTrend.description
    hide: @rollupMode.selected.mode != "direct"
    //animation: true
  // chart line #barChart {
  //   lineType: monotone
  //   lineWidth: 2
  //   dotSize: 5
  // }

    series {
      label: " "
      value: parseInt("a")
      chart bar {
        legendType: none
      }
    }
    series #user {
      label: @rollupMode.selectedLabel
      value: :dimensionScore()
      chart line {
        lineType: monotone
      }
    }


    scope filter {
      name: period
      value: AllPeriods
    }

    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }
    category cut #periods {
      value: .reportHistory:trendYear
      sortBy: .reportHistory:trendYear
      sortOrder: ascending
    }
    axis category {
      interval: preserveStartEnd
    }

    series #entire {
      label: "Overall Organization"
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      value: :dimensionScore()
      chart line {
        lineType: monotone
      }
    }

    series #benchmark {
      label: @defaultBenchmmark.selected.definitionName
      value: lookup value {
        source: benchmarks
        mapping value {
          value: @externalConfig.primaryDimensionId
          selector: bmValueCode
        }
        mapping value {
          value: @defaultBenchmmark.selected.definitionId
          selector: benchmarkDefinitionID
        }
        mapping header {
          header: periods
          selector: TrendYear
        }
        value: mean
        formatter: scoreFormatter
      }
      chart line {
        lineType: monotone
      }
      legend: rightMiddle
      axis primary {
      }
      axis secondary #secondaryAxis {
        hide: true
      }
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: medium
  } //here   
  widget headline #summaryDRLeaderIndex {
    label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
    description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
    hide: @rollupMode.selected.mode != "direct"

    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold." //what to display
    }
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVLeaderIndex.infoText
          label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: orgDetails
        }

      }
    }


    // suppressRule {
    //   criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected
    //   label: "The number of responses for your team is below the minimum threshold required to display results."
    // }

    cell: @dtEngagementSummary.m.data.main
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      //Area for labels
      area #labelFirst {
        width: '40%'
        display: block
        paddingLeft: 15px
      }
      // area #labelSecond {
      //   width: '30%'
      //   display: block
      //   //paddingLeft: 30px
      // }
      area #labelThird {
        display: block
        width: '50%'
        // paddingLeft: 10px
      }

      area #left {
        width: '35%'
        //display: block
        // height:300px
      }
      // area #middle {
      //   width: '30%'
      //   paddingLeft: 15px
      //   display: block
      //   height: 300px
      //   /* position: relative
      //   area #donut {
      //     position: absolute
      //   } */
      //   /* area #center {
      //     position: absolute
      //   } */
      // }
      area #right {
        width: '60%'
        display: block

      }
    }


    filter expression {
      value: .dimensions:id = "leaderindex"
    }

    //Text Tiles for Headers
    tile text #textTile_2 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelFirst
      value: "Overall Leader Index for Your Team"
    }
    // tile text #textTile_3 {
    //   style {
    //     fontSize: 16px
    //     fontWeight: bold
    //   }
    //   areaId: labelSecond
    //   value: "Group Distribution by Leader Index Score"
    // }
    tile text #textTile_4 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelThird
      value: "Items Included in Your Leader Index"
    }
    // tile text #textTile_5 {
    //   style {
    //     fontSize: 18px
    //     fontWeight: bold
    //   }
    //   areaId: labelThird
    //   value: "Mean Score"
    // }
    // tile text #textTile_6 {
    //   style {
    //     fontSize: 18px
    //     fontWeight: bold
    //   }
    //   areaId: labelFourth
    //   value: "Percentile Rank"
    // }

    //Chart and Table Tiles
    tile custom #leaderindex {

      areaId: left
      expression #score {
        value: :dimensionScore()//@cell.current
        valueFormatter: scoreFormatter
      }
      formula #change {
        value: @cell.change
        valueFormatter: scoreFormatter
      }
      expression #percentile {
        value: @dtEngagementSummary.m.data.benchmark.rank
        formatter: rankFormatter
      }
      expression #asteric {
        value: @cell.asteric//IIF(@cell.sig != 0, "*", " ")
      }
      expression #arrow {
        value: @cell.arrow//IIF(@cell.change > 0, "↑", IIF(change[] < 0, "↓", "-"))
      }
      expression #sigInfo {
        value: @cell.sigInfo// IIF(@cell.sig != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      formula #arrowColor {
        value: IIF(change[] > 0, IIF(@cell.sig != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(@cell.sig != 0, "#d02625", "Black"), "Black"))
      }
      formula #historyMean {
        value: @cell.current - @cell.change
        formatter: floatDefaultFormatter
      }
      // expression #score {
      //   value: :dimensionScore()
      //   valueFormatter: scoreFormatter
      // }
      expression #color {
        value: IIF(@cell.current >= 4, "#1FA583", IIF(@cell.current <= 2.5, "#D02525", "#E79F0B"))
      }
      expression #label {
        value: IIF(@cell.current >= 4, "High", IIF(@cell.current <= 2.5, "#D02525", "Moderate"))

      }
      //     formula #current {
      //       value: score[column = /history.current]
      //     }
      //     formula #change {
      //       value: diffSum[column = /history.current]
      //       formatter: floatDefaultFormatter
      //     }
      //     formula #arrow {
      //       //CNJ126 arrows ↑↓ or  ↑ ↓
      //       value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
      //     }
      //     formula #asteric {
      //       value: IIF(sig[column = /history.current] != 0, "*", " ")
      //     }
      formula #sigText {
        value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      //               formula #arrowColor {
      //       value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
      //     }
      //     formula #historyMean {
      //       value: score[column = /history.current] - diffSum[column = /history.current]
      //       formatter: floatDefaultFormatter
      //     }

      expression #description {
        value: IIF(:dimensionScore() >= 4, "Group is ready to have improvement planning discussions with their direct leader.", IIF(:dimensionScore() <= 2.5, "Focus should be placed on building relationships between direct leader and team prior to improvement planning.", "Group may be ready for improvement planning discussions, but the direct leader may benefit from additional guidance."))
      }
      //cb here

      formatString: '<span style= "margin-left:80px;font-size:60px"> {score}</span><span style ="color:{arrowColor}">{arrow}</span><br><span style="font-size:40px; margin-left:95px; color:{color};">{label}</span><br><br><p style="font-size:16px; margin-left:10px;">{description}</p>'
      // tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {arrowColor};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

    }
    // tile chartPlus #t1 {
    //   // filter expression {
    //   //   value: :combined_sourceid = "p494984785246"
    //   // }
    //   areaId: middle
    //   style {
    //     width: 500px
    //     height: 260px
    //     //paddingBottom: 10px
    //   }
    //   //test if palette work
    //   // palette: posNeuNeg

    //   axis primary #primaryAxis {
    //     hide: true
    //   }
    //   chartMargin {
    //     top: 40
    //   }
    //   series {
    //     label: "Responses"
    //     //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
    //     value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
    //     // removeEmptySeries: true
    //     base: count(unitHierarchy:)
    //     chart bar {
    //       // mode: stacked
    //       showBase: true
    //       valueLabel: "Groups"
    //       valuePosition: outer
    //     }
    //     format: percentNoDecimal
    //   }
    //   category cut {
    //     //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
    //     value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
    //     palette: LIpalette

    //   }
    // }




    tile grid #gridTile_2 {

      areaId: right
      style {
        width: "100%"
      }
      showBullets: false

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }

      row #headerLabels {
        label: " "
        cell custom {
          row: headerLabels
          column: main
          formula #value {
            value: "Mean Score"
          }
          formatString: "<b>{value}</b>"
        }
      }
      cell custom { //Errors out if you put too many cells 
        row: headerLabels
        column: benchmark
        formula #value {
          value: "Percentile Rank"
        }
        formatString: "<b>{value}</b>"
      }
      row list #items {
        table: .items:
        value: answerText(.items:Id) //toText(.items:SequenceId) + ". " + 
      }

      column cut #history {
        hide: true
        //categories: "'_1'"
        scope filter {
          name: period
          value: currentAndPrevious
        }
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :itemScore()
          }
          statistic mean #sig {
            testingType: T
            argument: numeric(.item_score:questionScoreValue)
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diffSum}"
          tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
        }
      }
      column #main {
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #asteric {
            value: IIF(sig[column = /history.current] != 0, "*", " ")
          }
          formula #sigText {
            value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
          }
          formula #historyMean {
            value: score[column = /history.current] - diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }

          formatString: "<pre>{current}<span style='color:{color};font-size:20px;'>{arrow}</span>{asteric}</pre>"
          tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        }
      }
      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: :itemScore()
            formatter: rankFormatter
          }
          lookup value #mean {
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: mean
            formatter: scoreFormatter
          }
          formula #tooltip {
            value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
            //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
          }
          formatString: "{rank}"
          tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
    //tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

        }
      }
    }
    size: medium
  }
  widget chart #summaryDRLeaderIndexChart {
    label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
    description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
    hide: @rollupMode.selected.mode != "direct"
    // st {
    // }
    filter expression {
      value: .dimensions:id = "leaderindex"
    }
    series #DRScore {
      label: "Your Score"
        //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
      value: :dimensionScore()
        // removeEmptySeries: true
        // base: count(unitHierarchy:)
      chart bar {
          // mode: stacked
          // showBase: true
          // valueLabel: "Groups"
        valuePosition: outer

      }
      format: scoreFormatter
    }
    series #OverallScore {
      label: "Organization"
      value: :dimensionScore()
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      chart bar {
          // mode: stacked
          // showBase: true
          // valueLabel: "Groups"
        valuePosition: outer

      }

    }

    axis category #categoryAxis {
    }
    axis primary #primaryAxis {

      format: percentNoDecimal
      minValue: 0
      maxValue: 5
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: medium
  }



  widget dataGrid #summaryDRKeyDrivers {
    label: @widgetConfig.lookup.data.summaryDRKeyDrivers.label
    description: @widgetConfig.lookup.data.summaryDRKeyDrivers.description
    size: medium
    hide: @rollupMode.selected.mode != "direct"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryDRKeyDrivers.infoText
          label: @widgetConfig.lookup.data.summaryDRKeyDrivers.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/score100"
      sortOrder: descending
      takeTop: 6
    }


   //filterexpression{ value: .dimension_score:dg1_dimensionScore = "Standard_3" }			

    row cut #itemsRow {
      total: none
      value: .item_score:dg1_questionScore
      //TODO: Need to exclude engagement items (filter out)
      // filter expression {
      //   value: .item_score:dg1_questionScore = "EV10137"      
      // }

    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:)
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint

        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }
    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }


    }



    column #gpr {
      label: "Percentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }

  widget dataGrid #summaryDRTopPerform {
    label: @widgetConfig.lookup.data.summaryDRTopPerform.label
    description: @widgetConfig.lookup.data.summaryDRTopPerform.description
    size: medium
    hide: @rollupMode.selected.mode != "direct"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryDRTopPerform.infoText
          label: @widgetConfig.lookup.data.summaryDRTopPerform.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/gpr"
      sortOrder: descending
      takeTop: 5
    }




   //filterexpression{ value: .dimension_score:dg1_dimensionScore = "Standard_3" }			

    row cut #itemsRow {
      total: none
      value: .item_score:dg1_questionScore
      //TODO: Need to exclude engagement items (filter out)
      // filter expression {
      //   value: .item_score:dg1_questionScore = "EV10137"      
      // }

    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:)
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint
        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }

    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }


    }



    column #gpr {
      label: "Precentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }

  widget dataGrid #summaryDRAddDimensions {
    label: @widgetConfig.lookup.data.summaryDRAddDimensions.label
    description: @widgetConfig.lookup.data.summaryDRAddDimensions.description
    hide: @rollupMode.selected.mode != "direct"
    size: large
    filter expression {
      value: .dimensions:includeHXWidget
    }
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryDRAddDimensions.infoText
          label: @widgetConfig.lookup.data.summaryDRAddDimensions.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }

    row list #dimensions {
      table: .dimensions:
      value: .dimensions:id
      total: none
    }

    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :dimensionScore()
        }
        statistic mean #sig {
          testingType: T
          argument: .dimension_score:dimensionScoreValue
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
      }
    }
    // column #recoding {
    //   label: " "
    //   cell custom {
    //     expression #type {
    //       value: ToText(.dimensions:id)
    //     }
    //     formula #teamIndex {
    //         //later should be recoce()
    //       value: IIF(value[column = /history.current] >= @externalConfig.teamIndex1, "TI-1", IIF(score[column = /history.current] < @externalConfig.teamIndex2, "TI-3", "TI-2"))
    //     }
    //     formula #team {
    //       value: IIF(type[] = "teamindex", teamIndex[])
    //     }

    //     formatString: "{team}"
    //   }
    // }
    column #main {
      label: "Mean score"
      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          //CNJ126 arrows ↑↓ or  ↑ ↓
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='font-size: 20px; color:{color};'>{arrow}</span>{asteric}</pre>"//To add Astric: 
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        // tooltipFormatString: "<b style='font-size:20px'>{historyMean}</b><br>Historical Mean Score" + "<br><b style='font-size:20px'>{change}</b><br> vs " + @surveyToCompareWith.selectedLabel + "<br><span style='  height: 25px;  width: 25px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }
    column #benchmark {
      label: "Percentile"
      cell custom {
        lookup rank #rank {
          takeInArray: Per
          mode percentile {
          }
          source: benchmarks
          mapping header {
            header: dimensions
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :dimensionScore()
          formatter: rankFormatter
        }
        lookup value #mean {
          source: benchmarks
          mapping header {
            header: dimensions
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: mean
          formatter: scoreFormatter
        }
        formula #tooltip {
          value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
        }
        formatString: "{rank}"
        tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>" + @defaultBenchmmark.selectedLabel + " Mean Score "
      }
    }
    column #recoding {
      label: " "
      sortable: false
      cell custom {
        formatString: " "
      }
    }

  }


}

page #Overall {

  label: "Overall"
  scope reportingHierarchy {
    reportingHierarchy: unitHierarchy
    mode: @rollupMode.selected.mode
  }
  dataTable #dtEngagementNodesOverall {
    dataGrid #dgEngagementNodesTMP {
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      scope filter {
        name: period
        value: currentAndPrevious
      }

      size: large
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }
      filter expression {
        value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
      }

      row list #nodes {
        total: none
        table: unitHierarchy:
        value: ""//unitHierarchy:language_text
        // takeTop: 5
        // sortBy: "/base"//count(:, .surveys:id = 1)
        take: 5
        sortBy: count(:, .reportHistory:historyTypeCode = "current")
        sortOrder: descending
      }

      column #nodeLabel {
        cell {
          value: unitHierarchy:language_text
        }
      }
      column #base {
        cell {
          value: count(:, .reportHistory:historyTypeCode = "current")
        }
      }
      column cut #history {
        // scope filter {
        //   name: period
        //   value: currentAndPrevious
        // }

        value: .reportHistory:historyTrendOrder
        total: none

        cell custom {
          expression #score {
            value: :dimensionScore()
          }
          statistic mean #sig {
            testingType: T
            argument: .dimension_score:dimensionScoreValue
            compare: next
          }

          formatString: "{score} [{sig}]"
        }
      }
      column #main { //This is where Engagement For your largest Groups is obtained from
        label: main
        cell custom {
          formula #score {
            value: score[column = /history.1]
          }
          formula #change {
            value: score[column = /history.1] - score[column = /history.2]
          }
          formula #sig {
            value: sig[column = /history.1]
          }
          formula #asteric {
            value: IIF(sig[] != 0, "*", " ")
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #historyMean {
            value: score[column = /history.2]
          }
          formula #sigInfo {
            value: IIF(sig[] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.1] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.1] != 0, "#d02625", "Black"), "Black"))
          }
          formatString: "{score} ({change}) [{sig}]"
        }
      }

      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarksById
            mapping value {
              value: @externalConfig.primaryDimensionId
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.idInt
              selector: BenchmarkId
            }
            value: :dimensionScore()
            formatter: rankFormatter
          }
          formatString: "{rank}"
        }
      }
      column #microchart {
        cell microchart {
          value: count(.dimension_score:)
          breakdownBy cut {
            value: .dimension_score:engagementFourPoint
          }
          microchart pie {
          }
        }
      }
    }
    map #m {
      from: nodes
    }
  }

  widget headline #overallResponseRate {
    label: @widgetConfig.lookup.data.overallResponseRate.label
    description: @widgetConfig.lookup.data.overallResponseRate.description
    size: large
    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    // Do not need to hide values on response rate widget
    // suppressRule {
    //   criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
    //   label: "Too few responses" //what to display
    // }
    // hide: @rollupMode.Selected.value

    toolbar { //start toolbar
      button #infobox {
        action showInfobox {
          info: @widgetConfig.lookup.data.overallResponseRate.infoText
          label: @widgetConfig.lookup.data.overallResponseRate.label
          size: large
        }
      }
      button #export {
        action export {
          format: png
        }
      }
      button #navigate {
        action navigate {
          navigateTo: response_rates
        }
      }
    } //end toolbar
    container: container flex {
      flexDirection: row
      flexWrap: wrap

      area #area_one_space {
        width: '7%'
        display: block
      }
      area #area_one {
        width: '9%'
        display: block
        verticalAlign: "center"
      }
      area #area_two {
        width: '13%'
        display: block
      }
      area #area_three_space {
        width: '12%'
        display: block
      }
      area #area_three {
        width: '5%'
        display: block
      }
      area #area_four {
        width: '14%'
        display: block
      }
      area #area_five_space {
        width: '11%'
        display: block
      }
      area #area_five {
        width: '5%'
        display: block
      }
      area #area_six {
        width: '16%'
        display: block
      }
    }
    tile text #textTile_01 {
      areaId: area_two
      value: "Response Rate"
      style {
        fontSize: 24
      }

    }

    tile value #valueTile_1 {
      areaId: area_two
      value: 100 * @cp.WFComplete / COUNT(:responseid)
      valueFormatter: percentNoDecimal
      style {
        fontSize: 40
        //fontWeight: bold
        color: #000000
        A {
        }

      }
      valueColorFormatter: dropOffDefaultFormatter
    }
    tile chartPlus #icon1 {
      areaId: area_one
      palette: icon_pie_palette
      style {
        height: 100px
      }
      chart pie {
        innerRadius: 30
        outerRadius: 45
        legendType: circle
      }
      series {
        label: "Responses"
        value: COUNT(:responseid) / count(:, true, "__top") * 100
        base: COUNT(:responseid)
        valueFormatter: statisticPercentsDefaultFormatter
      }
      category cut {
        value: :status
      }
      removeEmptyCategories: true


    }
    tile text #textTile_02 {
      areaId: area_four
      value: "Number Invited"
      style {
        fontSize: 24
        color: #000000
      }
    }
    tile value #valueTile_4 {
      areaId: area_four
      value: COUNT(:responseid)
      valueFormatter: bigNumberFormatter
      style {
        fontSize: 40
        color: #000000
      }
    }
    tile text #textTile_03 {
      areaId: area_six
      value: "Completed Surveys"
      style {
        fontSize: 24
      }
    }
    tile value #valueTile_3 {
      areaId: area_six
      value: @cp.WFComplete
      valueFormatter: bigNumberFormatter
      style {
        fontSize: 40
        color: #000000

      }
    }
    tile image #imageTile {
      areaId: area_three
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/file%20library%20test/RR_Invite.jpg"
    }
    tile image #imageTile_2 {
      areaId: area_five
      value: "/isa/BDJPFRDMEYBPBKLVADAYFQCDAVIOEQJR/file%20library%20test/RR_Complete.jpg"
    }
  }

  widget headline #overallPrimaryDimDonut {
    label: @widgetConfig.lookup.data.overallPrimaryDimDonut.label
    description: @widgetConfig.lookup.data.overallPrimaryDimDonut.description
  // hide: @rollupMode.selected.mode != "rollup"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.overallPrimaryDimDonut.infoText
          label: @widgetConfig.lookup.data.overallPrimaryDimDonut.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {
        action navigate {
          navigateTo: orgDetails
        }
      }
    }

    cell: @dtEngagementSummary.m.data.main
    //CNJ126 replaced container
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      area #labelFirst {
        width: '29%'
        display: block
        paddingLeft: 15px
      }
      area #labelSecond {
        display: block
        width: '60%'
        paddingLeft: 60px
      }
      // area #labelThird {
      //   display: block
      //   width: '35%'
      //   paddingLeft: 30px
      // }
      area #left {
        width: '30%'
        height: 300px
        paddingLeft: 50px

        position: relative
        area #donut {
          position: absolute
        }
        area #center {
          position: absolute
        }
      }
      // area #legend {
      //   width: '15%'
      //   display: flex
      //   flexDirection: column
      //   alignItems: baseline
      // }


      area #right {
        width: '70%'
        display: block
        paddingLeft: 30px
        paddingBottom: 30px
      }
      area #legend {
        width: '100%'
        paddingLeft: 20px
        paddingBottom: 30px

      }
    }


    filter expression {
      value: .dimensions:id = "engagement"
    }
    tile text #textTile_3 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelFirst
      value: "Engagement Mean Score and Level Distribution"
    }
    tile text #textTile_4 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelSecond
      value: "Items Included in Your Engagement Score"

    }
    // tile text #textTile_5 {
    //   style {
    //     fontSize: 16px
    //     fontWeight: bold
    //   }
    //   areaId: labelThird
    //   value: "Items Included in Your Engagement Score"
    // }

    tile microchart #microchartTile_2 {
      areaId: donut
      value: @dtEngagementSummary.m.data.microchart.value
      microchart pie {
        donutWidth: 30%
        percentFormat: percentNoDecimal
        //CNJ126 legend
        legendType: diamond
        palette: engaged
      }
      style {
        width: "350px"
        height: "250px"
      }
      legend: bottomCenter

    }


    tile custom #customTile_2 {
      areaId: center
      expression #score {
        value: @cell.current
        valueFormatter: scoreFormatter
      }
      expression #change {
        value: @cell.change
        valueFormatter: scoreFormatter
      }
      expression #percentile {
        value: @dtEngagementSummary.m.data.benchmark.rank
        formatter: rankFormatter
      }
      expression #asteric {
        value: @cell.asteric//IIF(@cell.sig != 0, "*", " ")
      }
      expression #arrow {
        value: @cell.arrow//IIF(@cell.change > 0, "↑", IIF(change[] < 0, "↓", "-"))
      }
      expression #sigInfo {
        value: @cell.sigInfo// IIF(@cell.sig != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      formula #color {
        value: IIF(change[] > 0, IIF(@cell.sig != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(@cell.sig != 0, "#d02625", "Black"), "Black"))
      }
      formula #historyMean {
        value: @cell.current - @cell.change
        formatter: floatDefaultFormatter
      }
      //CNJ126 arrows edited formatstring
      formatString: '{score} <span style="color:{color}">{arrow}</span> {asteric}<span style="font-size: 16px; color:grey; display:block">{percentile} percentile</span>'
      tooltipFormatString: "<span style='font-size:40px'>{historyMean}</span><br>Mean Score for " + @surveyToCompareWith.selectedLabel + "<br><br><span style='font-size:30px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigInfo}"

      style {
        fontSize: 40px
        display: block
        textAlign: center
      }
    }

    //CNJ126 Tile legend  For different legends; try ● ■
     //but then you should also change legendtype on Key drivers, datagrids and tooltips
    tile custom #legend_1 {
      areaId: legend
      formatString: '<span style="color:#027580"> ✦ </span> Highly Engaged'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_2 {
      areaId: legend
      formatString: '<span style="color:#1BA583">✦ </span> Engaged'
      style {
        fontSize: 14
      }
    }
    tile custom #legend_3 {
      areaId: legend
      formatString: '<span style="color:#E69F0D">✦ </span> Neutral'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_4 {
      areaId: legend
      formatString: '<span style="color:#D02624">✦ </span> Disengaged'
      style {
        fontSize: 14
      }
    }

    // tile chartPlus #summaryMTVTrend {
    //   label: @widgetConfig.lookup.data.summaryMTVTrend.label
    //   description: @widgetConfig.lookup.data.summaryMTVTrend.description
    //   hide: @rollupMode.selected.mode != "rollup"
    //   areaId: middle

    //   scope filter {
    //     name: period
    //     value: AllPeriods
    //   }


    //   filter expression {
    //     value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    //   }
    //   category cut #periods {
    //     value: .reportHistory:trendYear
    //     sortBy: .reportHistory:trendYear
    //     sortOrder: ascending
    //   }

    //   series {
    //     label: ""
    //     value: parseInt("a")
    //     chart bar {
    //       legendType: none
    //     }
    //   }

    //   axis category {
    //     interval: preserveStartEnd
    //   }

    //   series #user {
    //     label: @rollupMode.selectedLabel
    //     value: :dimensionScore()
    //     chart line {
    //     }
    //   }
    //   series #entire {
    //     label: "Entire organization"
    //     scope reportingHierarchy {
    //       reportingHierarchy: unitHierarchy
    //       nodes: AllData
    //     }
    //     filter expression {
    //       value: _isNotNull(@unitHierarchy.source)
    //     }
    //     value: :dimensionScore()
    //     chart line {
    //     }
    //   }
    //   series #benchm {

    //     label: @defaultBenchmmark.selected.definitionName
    //     value: lookup value {
    //       source: benchmarks
    //       mapping value {
    //         value: @externalConfig.primaryDimensionId
    //         selector: bmValueCode
    //       }
    //       mapping value {
    //         value: @defaultBenchmmark.selected.definitionId
    //         selector: benchmarkDefinitionID
    //       }
    //       mapping header {
    //         header: periods
    //       //value: .reportHistory:trendYear
    //         selector: TrendYear
    //       }
    //       value: mean
    //       formatter: scoreFormatter
    //     }
    //     chart line {
    //     }
    //   }
    //   legend: rightMiddle
    //   axis primary {
    //   }

    //   axis secondary #secondaryAxis {
    //     hide: true
    //   }
    // }


    tile grid #gridTile_2 {

      areaId: right
      style {
        width: "100%"
      }
      showBullets: false

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }
      row #headerLabels {
        label: " "
        cell custom {
          row: headerLabels
          column: main
          formula #value {
            value: "Mean Score"
          }
          formatString: "<b>{value}</b>"
        }
      }
      cell custom { //Errors out if you put too many cells 
        row: headerLabels
        column: benchmark
        formula #value {
          value: "Percentile Rank"
        }
        formatString: "<b>{value}</b>"
      }
      row list #items {
        table: .items:
        value: answerText(.items:Id) //toText(.items:SequenceId) + ". " +
      }

      column cut #history {
        hide: true
        //categories: "'_1'"
        scope filter {
          name: period
          value: currentAndPrevious
        }
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :itemScore()
          }
          statistic mean #sig {
            testingType: T
            argument: numeric(.item_score:questionScoreValue)
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diffSum}"
          tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

        }
      }
      column #main {
        label: "Mean Score"
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #asteric {
            value: IIF(sig[column = /history.current] != 0, "*", " ")
          }
          formula #sigText {
            value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.1] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
          }
          formula #historyMean {
            value: score[column = /history.current] - diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }

          formatString: "<pre>{current}<span style='font-size:20px; color:{color};'>{arrow}</span>{asteric}</pre>"
          tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        }
      }
      column #benchmark {
        cell custom {
          lookup rank #rank {

            takeInArray: Per
            mode percentile {
              ends: tonearest
            }
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: :itemScore()
            formatter: rankFormatter
          }
          lookup value #mean {
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: mean
            formatter: scoreFormatter
          }
          formula #tooltip {
            value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>Benchmark Mean Value: " + mean[], "too few responses")
            //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
          }
          formatString: "{rank}"
          tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
    //          tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

        }
      }
    }
    size: halfwidth
  }
  widget chart #overallTrend {
    label: @widgetConfig.lookup.data.overallTrend.label
    description: @widgetConfig.lookup.data.overallTrend.description
  // hide: @rollupMode.selected.mode != "rollup"
    //animation: true
  // chart line #barChart {
  //   lineType: monotone
  //   lineWidth: 2
  //   dotSize: 5
  // }
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    series {
      label: " "
      value: parseInt("a")
      chart bar {
        legendType: none
      }
    }
    series #user {
      label: @rollupMode.selectedLabel
      value: :dimensionScore()
      chart line {
        lineType: monotone
      }
    }


    scope filter {
      name: period
      value: AllPeriods
    }

    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }
    category cut #periods {
      value: .reportHistory:trendYear
      sortBy: .reportHistory:trendYear
      sortOrder: ascending
    }
    axis category {
      interval: preserveStartEnd
    }

    series #entire {
      label: "Overall Organization"
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      value: :dimensionScore()
      chart line {
        lineType: monotone
      }
    }

    series #benchmark {
      label: @defaultBenchmmark.selected.definitionName
      value: lookup value {
        source: benchmarks
        mapping value {
          value: @externalConfig.primaryDimensionId
          selector: bmValueCode
        }
        mapping value {
          value: @defaultBenchmmark.selected.definitionId
          selector: benchmarkDefinitionID
        }
        mapping header {
          header: periods
          selector: TrendYear
        }
        value: mean
        formatter: scoreFormatter
      }
      chart line {
        lineType: monotone
      }
      legend: rightMiddle
      axis primary {
      }
      axis secondary #secondaryAxis {
        hide: true
      }
    }
    axis primary #primaryAxis {
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: medium
  } //here   
  widget headline #overallLargeGroups {

    size: large
    label: @widgetConfig.lookup.data.overallLargeGroups.label
    description: @widgetConfig.lookup.data.overallLargeGroups.description
    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected
      label: "The number of responses for your team is below the minimum theshold required to display results."
    }
    toolbar {
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.overallLargeGroups.infoText
          label: @widgetConfig.lookup.data.overallLargeGroups.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }
      button #navigate {
        action navigate {
          navigateTo: page_5
        }
          // action setSelector {
          //   value: Engagement
          //    select: @dimensionsSelector2
          // }
      }
    }

    //CNJ126 padding botttom
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      area #donuts {
        width: '100%'
        display: flex
        paddingLeft: 30px
        paddingBottom: 30px
        justifyContent: "center"//"space-evenly"
      }
      area #legend {
        width: '100%'
        paddingLeft: 20px
        paddingBottom: 30px

      }
    }


    tile set #setTile_2 {
      areaId: donuts
      //CNJ126 tileset switch container flex with grid
      container: container grid {
        rows: 'A A A A A'
        justifyContent: spaceEvenly

      }
      /* container: container flex {
        flexDirection: row
        flexWrap: wrap
      } */

      itemContainer: container flex {
        flexDirection: column
          // backgroundColor: yellow
        width: 300px
          //display: flex

        area #label {
          height: 50px
          display: block
        }
        area #respondents {
            // height: 10px
          display: block
        }
        area #main {
          //  width: 500px
          //  height: 500px
            // backgroundColor: orange
          position: relative
          area #donut {
              // backgroundColor: green
              //position: absolute
              // top: "50%"
              // left: "50%"
              // transform: "translate(-50%, -50%)"
          }
          area #center {
              // backgroundColor: orange
            position: absolute
              // top: "50%"
              // left: "50%"
              // transform: "translate(-50%, -50%)"
          }
        }
      }

      breakdownBy inlineData {
        value: @dtEngagementNodesOverall.m.data
      }

      tile text {
        areaId: label
        value: this.nodeLabel.value
        style {
          fontSize: 15px
          //fontWeight: bold
        }
      }
      tile value {
        areaId: respondents
        value: this.base.value
        formatString: "{value} Responses"
        style {
          fontSize: 16px
        }
      }

      tile microchart {
        areaId: donut
        value: this.microchart.value

        microchart pie {
          donutWidth: 30px
          palette: engaged
          valuePosition: outer
          percentFormat: percentNoDecimal

        }
        style {
          height: 205px
          width: 260px
            // paddingBottom:25px

        }
      }


      tile custom #customTile_2 {
        areaId: center
        expression #score {
          value: this.main.score
          valueFormatter: scoreFormatter
        }
        expression #change {
          value: this.main.change
          valueFormatter: scoreFormatter
        }
        expression #percentile {
          value: this.benchmark.rank
          formatter: rankFormatter
        }
        expression #asteric {
          value: this.main.asteric//IIF(this.main.sig != 0, "*", " ")
        }
        expression #arrow {
          value: this.main.arrow//IIF(this.main.change > 0, "↑", IIF(this.main.change < 0, "↓", "-"))
        }
        expression #sigInfo {
          value: this.main.sigInfo//IIF(this.main.sig != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        expression #label {
          value: this.main.label
        }
        expression #color {
          value: this.main.color
        }
        expression #historyMean {
          value: this.main.historyMean
        }
      //CNJ126 arrows edited formatstring
        formatString: '<span style="font-size: 30px; display:block">{score} <span style="color:{color}">{arrow}</span> {asteric}</span><span style="font-size: 14px; color:grey; display:block">{percentile} Percentile</span>'
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigInfo}"


          // formatString: '{score} {arrow} {asteric}<span style="font-size: 20px; display:block">{percentile} percentile</span>'
          // tooltipFormatString: "change {change} vs {}label}" + "<br/>{sigInfo}"

        style {
          fontSize: 40px
          display: block
          textAlign: center
        }
      }



    }

    tile custom #legend_1 {
      areaId: legend
      formatString: '<span style="color:#027580"> ✦ </span> Highly Engaged'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_2 {
      areaId: legend
      formatString: '<span style="color:#1BA583">✦ </span> Engaged'
      style {
        fontSize: 14
      }
    }
    tile custom #legend_3 {
      areaId: legend
      formatString: '<span style="color:#E69F0D">✦ </span> Neutral'
      style {
        fontSize: 14
      }
    }

    tile custom #legend_4 {
      areaId: legend
      formatString: '<span style="color:#D02624">✦ </span> Disengaged'
      style {
        fontSize: 14
      }
    }

  }

  // widget headline #summaryMTVLeaderIndex {
  //   label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
  //   description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
  //   hide: @rollupMode.selected.mode != "rollup"

  //   suppressRule {
  //     criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected //when
  //     label: "The number of responses for your team is below the minimum threshold." //what to display
  //   }
  //   toolbar { // This 
  //     button #infobox {
  //       action showInfobox {
  //         size: large
  //         info: @widgetConfig.lookup.data.summaryMTVLeaderIndex.infoText
  //         label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
  //       }
  //     }
  //     button #export {
  //       action export {
  //         format: png
  //       }
  //     }

  //     button #navigate {

  //       action navigate {
  //         navigateTo: orgDetails
  //       }

  //     }
  //   }


  //   // suppressRule {
  //   //   criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected
  //   //   label: "The number of responses for your team is below the minimum threshold required to display results."
  //   // }

  //   cell: @dtEngagementSummary.m.data.main
  //   container: container flex {
  //     flexDirection: row
  //     flexWrap: wrap
  //     //Area for labels
  //     area #labelFirst {
  //       width: '29%'
  //       display: block
  //       paddingLeft: 40px
  //       // paddingBottom:20px
  //     }
  //     area #labelSecond {
  //       width: '30%'
  //       display: block
  //       paddingLeft: 30px
  //     }
  //     area #labelThird {
  //       display: block
  //       width: '40%'

  //     }
  //     // area #labelFourth {
  //     //   display: block
  //     //   width: '7%'
  //     //   // paddingLeft: 34px
  //     // }
  //     //Area for charts and tables
  //     area #left {
  //       width: "25%"
  //     }
  //     area #middle {
  //       width: "30%"
  //       paddingLeft: 40px
  //       height: 400px
  //       position: relative
  //       area #donut {
  //         position: absolute
  //       }
  //       area #center {
  //         position: absolute
  //       }
  //     }
  //     area #right {
  //       width: "40%"
  //       //paddingLeft: 40px
  //     }
  //   }


  //   filter expression {
  //     value: .dimensions:id = "leaderindex"
  //   }

  //   //Text Tiles for Headers
  //   tile text #textTile_2 {
  //     style {
  //       fontSize: 16px
  //       fontWeight: bold
  //     }
  //     areaId: labelFirst
  //     value: "Overall Leader Index for Your Team"
  //   }
  //   tile text #textTile_3 {
  //     style {
  //       fontSize: 16px
  //       fontWeight: bold
  //     }
  //     areaId: labelSecond
  //     value: "Group Distribution by Leader Index Score"
  //   }
  //   tile text #textTile_4 {
  //     style {
  //       fontSize: 16px
  //       fontWeight: bold
  //     }
  //     areaId: labelThird
  //     value: "Items Included in Your Leader Index"
  //   }
  //   // tile text #textTile_5 {
  //   //   style {
  //   //     fontSize: 18px
  //   //     fontWeight: bold
  //   //   }
  //   //   areaId: labelThird
  //   //   value: "Mean Score"
  //   // }
  //   // tile text #textTile_6 {
  //   //   style {
  //   //     fontSize: 18px
  //   //     fontWeight: bold
  //   //   }
  //   //   areaId: labelFourth
  //   //   value: "Percentile Rank"
  //   // }

  //   //Chart and Table Tiles
  //   tile custom #leaderindex {
  //     expression #score {
  //       value: :dimensionScore()
  //       valueFormatter: scoreFormatter
  //     }
  //     expression #color {
  //       value: IIF(:dimensionScore() >= 4, "#1FA583", IIF(:dimensionScore() <= 2.5, "#D02525", "#E79F0B"))
  //     }
  //     expression #label {
  //       value: IIF(:dimensionScore() >= 4, "High", IIF(:dimensionScore() <= 2.5, "#D02525", "Moderate"))

  //     }
  //     expression #description {
  //       value: IIF(:dimensionScore() >= 4, "Group is ready to have improvement planning discussions with their direct leader.", IIF(:dimensionScore() <= 2.5, "Focus should be placed on building relationships between direct leader and team prior to improvement planning.", "Group may be ready for improvement planning discussions, but the direct leader may benefit from additional guidance."))
  //     }
  //   //cb here
  //     areaId: left

  //     formatString: '<span style= "margin-left:200px;"><span style="font-size:60px";> {score}</span><br><span style="font-size:40px; margin-left:210px; color:{color};">{label}</span><br><br><p style="font-size:16px; margin-left:30px;">{description}</p>'

  //   }
  //   tile chartPlus #t1 {
  //     // filter expression {
  //     //   value: :combined_sourceid = "p494984785246"
  //     // }
  //     areaId: donut
  //     style {
  //       width: 350px
  //       paddingBottom: 10px
  //     }
  //     //test if palette work
  //     // palette: posNeuNeg

  //     axis primary #primaryAxis {
  //       hide: true
  //     }
  //     chartMargin {
  //       top: 40
  //     }
  //     series {
  //       label: "Responses"
  //       //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
  //       value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
  //       // removeEmptySeries: true
  //       base: count(unitHierarchy:)
  //       chart bar {
  //         // mode: stacked
  //         showBase: true
  //         valueLabel: "Groups"
  //         valuePosition: outer
  //       }
  //       format: percentNoDecimal
  //     }
  //     category cut {
  //       //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
  //       value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
  //       palette: LIpalette

  //     }
  //   }




  //   tile grid #gridTile_2 {

  //     areaId: right
  //     style {
  //       width: "100%"
  //     }
  //     showBullets: false

  //     suppression recordsBase {
  //       threshold: @suppressionThreshold.selected
  //     }

  //     row #headerLabels {
  //       label: " "
  //       cell custom {
  //         row: headerLabels
  //         column: main
  //         formula #value {
  //           value: "Mean Score"
  //         }
  //         formatString: "<b>{value}</b>"
  //       }
  //     }
  //     cell custom { //Errors out if you put too many cells 
  //       row: headerLabels
  //       column: benchmark
  //       formula #value {
  //         value: "Percentile Rank"
  //       }
  //       formatString: "<b>{value}</b>"
  //     }
  //     row list #items {
  //       table: .items:
  //       value: answerText(.items:Id) //toText(.items:SequenceId) + ". " + 
  //     }

  //     column cut #history {
  //       hide: true
  //       //categories: "'_1'"
  //       scope filter {
  //         name: period
  //         value: currentAndPrevious
  //       }
  //       total: none
  //       value: .reportHistory:historyTypeCode
  //       cell custom {
  //         expression #score {
  //           value: :itemScore()
  //         }
  //         statistic mean #sig {
  //           testingType: T
  //           argument: numeric(.item_score:questionScoreValue)
  //           compare: next
  //         }
  //         formula #diff {
  //           value: score[column = %.current] - score[]
  //         }
  //         formula #diffSum {
  //           value: sum(diff[column = %.*])
  //         }
  //         formatString: "{score} [{sig}] {diffSum}"
  //         tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
  //       }
  //     }
  //     column #main {
  //       cell custom {
  //         formula #current {
  //           value: score[column = /history.current]
  //         }
  //         formula #change {
  //           value: diffSum[column = /history.current]
  //           formatter: floatDefaultFormatter
  //         }
  //         formula #arrow {
  //           //CNJ126 arrows ↑↓ or  ↑ ↓
  //           value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
  //         }
  //         formula #asteric {
  //           value: IIF(sig[column = /history.current] != 0, "*", " ")
  //         }
  //         formula #sigText {
  //           value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
  //         }
  //         formula #color {
  //           value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
  //         }
  //         formula #historyMean {
  //           value: score[column = /history.current] - diffSum[column = /history.current]
  //           formatter: floatDefaultFormatter
  //         }
  //         formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
  //         tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

  //       }
  //     }
  //     column #benchmark {
  //       cell custom {
  //         lookup rank #rank {
  //           takeInArray: Per
  //           mode percentile {
  //           }
  //           source: benchmarks
  //           mapping header {
  //             header: items
  //             selector: bmValueCode
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.definitionId
  //             selector: BenchmarkDefinitionId
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.periodId
  //             selector: TrendYear
  //           }
  //           value: :itemScore()
  //           formatter: rankFormatter
  //         }
  //         lookup value #mean {
  //           source: benchmarks
  //           mapping header {
  //             header: items
  //             selector: bmValueCode
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.definitionId
  //             selector: BenchmarkDefinitionId
  //           }
  //           mapping value {
  //             value: @defaultBenchmmark.selected.periodId
  //             selector: TrendYear
  //           }
  //           value: mean
  //           formatter: scoreFormatter
  //         }
  //         formula #tooltip {
  //           value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
  //           //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
  //         }
  //         formatString: "{rank}"
  //         tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
  //   //tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

  //       }
  //     }
  //   }
  //   size: large
  // }

  widget headline #overallLeaderIndex {
    label: @widgetConfig.lookup.data.overallLeaderIndex.label
    description: @widgetConfig.lookup.data.overallLeaderIndex.description
  // hide: @rollupMode.selected.mode != "rollup"
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold." //what to display
    }
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.overallLeaderIndex.infoText
          label: @widgetConfig.lookup.data.overallLeaderIndex.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: orgDetails
        }

      }
    }


    // suppressRule {
    //   criteria: count(:, .reportHistory:id = 1001) < @suppressionThreshold.selected
    //   label: "The number of responses for your team is below the minimum threshold required to display results."
    // }

    cell: @dtEngagementSummary.m.data.main
    container: container flex {
      flexDirection: row
      flexWrap: wrap
      //Area for labels
      area #labelFirst {
        width: '40%'
        display: block
        paddingLeft: 15px
      }
      // area #labelSecond {
      //   width: '30%'
      //   display: block
      //   //paddingLeft: 30px
      // }
      area #labelThird {
        display: block
        width: '50%'
        // paddingLeft: 10px
      }

      area #left {
        width: '35%'
        //display: block
        // height:300px
      }
      // area #middle {
      //   width: '30%'
      //   paddingLeft: 15px
      //   display: block
      //   height: 300px
      //   /* position: relative
      //   area #donut {
      //     position: absolute
      //   } */
      //   /* area #center {
      //     position: absolute
      //   } */
      // }
      area #right {
        width: '60%'
        display: block

      }
    }


    filter expression {
      value: .dimensions:id = "leaderindex"
    }

    //Text Tiles for Headers
    tile text #textTile_2 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelFirst
      value: "Overall Leader Index for Your Team"
    }
    // tile text #textTile_3 {
    //   style {
    //     fontSize: 16px
    //     fontWeight: bold
    //   }
    //   areaId: labelSecond
    //   value: "Group Distribution by Leader Index Score"
    // }
    tile text #textTile_4 {
      style {
        fontSize: 16px
        fontWeight: bold
      }
      areaId: labelThird
      value: "Items Included in Your Leader Index"
    }
    // tile text #textTile_5 {
    //   style {
    //     fontSize: 18px
    //     fontWeight: bold
    //   }
    //   areaId: labelThird
    //   value: "Mean Score"
    // }
    // tile text #textTile_6 {
    //   style {
    //     fontSize: 18px
    //     fontWeight: bold
    //   }
    //   areaId: labelFourth
    //   value: "Percentile Rank"
    // }

    //Chart and Table Tiles
    tile custom #leaderindex {

      areaId: left
      expression #score {
        value: @cell.current
        valueFormatter: scoreFormatter
      }
      expression #change {
        value: @cell.change
        valueFormatter: scoreFormatter
      }
      expression #percentile {
        value: @dtEngagementSummary.m.data.benchmark.rank
        formatter: rankFormatter
      }
      expression #asteric {
        value: @cell.asteric//IIF(@cell.sig != 0, "*", " ")
      }
      expression #arrow {
        value: @cell.arrow//IIF(@cell.change > 0, "↑", IIF(change[] < 0, "↓", "-"))
      }
      expression #sigInfo {
        value: @cell.sigInfo// IIF(@cell.sig != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      formula #arrowColor {
        value: IIF(change[] > 0, IIF(@cell.sig != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(@cell.sig != 0, "#d02625", "Black"), "Black"))
      }
      formula #historyMean {
        value: @cell.current - @cell.change
        formatter: floatDefaultFormatter
      }
      // expression #score {
      //   value: :dimensionScore()
      //   valueFormatter: scoreFormatter
      // }
      expression #color {
        value: IIF(@cell.current >= 4, "#1FA583", IIF(@cell.current <= 2.5, "#D02525", "#E79F0B"))
      }
      expression #label {
        value: IIF(@cell.current >= 4, "High", IIF(@cell.current <= 2.5, "#D02525", "Moderate"))

      }
      //     formula #current {
      //       value: score[column = /history.current]
      //     }
      //     formula #change {
      //       value: diffSum[column = /history.current]
      //       formatter: floatDefaultFormatter
      //     }
      //     formula #arrow {
      //       //CNJ126 arrows ↑↓ or  ↑ ↓
      //       value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
      //     }
      //     formula #asteric {
      //       value: IIF(sig[column = /history.current] != 0, "*", " ")
      //     }
      formula #sigText {
        value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
      }
      //               formula #arrowColor {
      //       value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
      //     }
      //     formula #historyMean {
      //       value: score[column = /history.current] - diffSum[column = /history.current]
      //       formatter: floatDefaultFormatter
      //     }

      expression #description {
        value: IIF(:dimensionScore() >= 4, "Group is ready to have improvement planning discussions with their direct leader.", IIF(:dimensionScore() <= 2.5, "Focus should be placed on building relationships between direct leader and team prior to improvement planning.", "Group may be ready for improvement planning discussions, but the direct leader may benefit from additional guidance."))
      }
      //cb here

      formatString: '<span style= "margin-left:80px;font-size:60px"> {score}</span><span style ="color:{arrowColor}">{arrow}</span><br><span style="font-size:40px; margin-left:95px; color:{color};">{label}</span><br><br><p style="font-size:16px; margin-left:10px;">{description}</p>'
      // tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {arrowColor};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

    }
    // tile chartPlus #t1 {
    //   // filter expression {
    //   //   value: :combined_sourceid = "p494984785246"
    //   // }
    //   areaId: middle
    //   style {
    //     width: 500px
    //     height: 260px
    //     //paddingBottom: 10px
    //   }
    //   //test if palette work
    //   // palette: posNeuNeg

    //   axis primary #primaryAxis {
    //     hide: true
    //   }
    //   chartMargin {
    //     top: 40
    //   }
    //   series {
    //     label: "Responses"
    //     //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
    //     value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
    //     // removeEmptySeries: true
    //     base: count(unitHierarchy:)
    //     chart bar {
    //       // mode: stacked
    //       showBase: true
    //       valueLabel: "Groups"
    //       valuePosition: outer
    //     }
    //     format: percentNoDecimal
    //   }
    //   category cut {
    //     //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
    //     value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
    //     palette: LIpalette

    //   }
    // }




    tile grid #gridTile_2 {

      areaId: right
      style {
        width: "100%"
      }
      showBullets: false

      suppression recordsBase {
        threshold: @suppressionThreshold.selected
      }

      row #headerLabels {
        label: " "
        cell custom {
          row: headerLabels
          column: main
          formula #value {
            value: "Mean Score"
          }
          formatString: "<b>{value}</b>"
        }
      }
      cell custom { //Errors out if you put too many cells 
        row: headerLabels
        column: benchmark
        formula #value {
          value: "Percentile Rank"
        }
        formatString: "<b>{value}</b>"
      }
      row list #items {
        table: .items:
        value: answerText(.items:Id) //toText(.items:SequenceId) + ". " + 
      }

      column cut #history {
        hide: true
        //categories: "'_1'"
        scope filter {
          name: period
          value: currentAndPrevious
        }
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :itemScore()
          }
          statistic mean #sig {
            testingType: T
            argument: numeric(.item_score:questionScoreValue)
            compare: next
          }
          formula #diff {
            value: score[column = %.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = %.*])
          }
          formatString: "{score} [{sig}] {diffSum}"
          tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
        }
      }
      column #main {
        cell custom {
          formula #current {
            value: score[column = /history.current]
          }
          formula #change {
            value: diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }
          formula #arrow {
            //CNJ126 arrows ↑↓ or  ↑ ↓
            value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
          }
          formula #asteric {
            value: IIF(sig[column = /history.current] != 0, "*", " ")
          }
          formula #sigText {
            value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
          }
          formula #color {
            value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
          }
          formula #historyMean {
            value: score[column = /history.current] - diffSum[column = /history.current]
            formatter: floatDefaultFormatter
          }

          formatString: "<pre>{current}<span style='color:{color};font-size:20px;'>{arrow}</span>{asteric}</pre>"
          tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        }
      }
      column #benchmark {
        cell custom {
          lookup rank #rank {
            takeInArray: Per
            mode percentile {
            }
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: :itemScore()
            formatter: rankFormatter
          }
          lookup value #mean {
            source: benchmarks
            mapping header {
              header: items
              selector: bmValueCode
            }
            mapping value {
              value: @defaultBenchmmark.selected.definitionId
              selector: BenchmarkDefinitionId
            }
            mapping value {
              value: @defaultBenchmmark.selected.periodId
              selector: TrendYear
            }
            value: mean
            formatter: scoreFormatter
          }
          formula #tooltip {
            value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
            //"<pre>" + current[] + " " + arrow[] + " " + asteric[] + "</pre>", "too few responses" )
          }
          formatString: "{rank}"
          tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>Benchmark Mean Value "
    //tooltipFormatString: "{tooltip}"//"percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value {mean}"

        }
      }
    }
    size: medium
  }

  widget chart #summaryMTVLeaderIndexChart {
    label: @widgetConfig.lookup.data.summaryMTVLeaderIndex.label
    description: @widgetConfig.lookup.data.summaryMTVLeaderIndex.description
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }
    series {
      label: "Responses"
        //value: count(:) / count(:, some(.dimension_score:, true, :), "__top") * 100
      value: count(unitHierarchy:) / count(unitHierarchy:, some(.dimension_score:, true, unitHierarchy:), "__top") * 100
        // removeEmptySeries: true
      base: count(unitHierarchy:)
      chart bar {
          // mode: stacked
        showBase: true
        valueLabel: "Groups"
        valuePosition: outer
        maxBarSize: 125

      }
      format: percentNoDecimal
    }
    category cut {
        //value: recode(avg(.dimension_score:dimensionScoreValue , true, :), @LeaderIndexGroup)
      value: recode(avg(.dimension_score:dimensionScoreValue, true, unitHierarchy:), @LeaderIndexGroup)
      palette: LIpalette

    }
    axis category #categoryAxis {
    }
    axis primary #primaryAxis {

      format: percentNoDecimal
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    size: medium
  }


  widget dataGrid #overallKeyDrivers {
    label: @widgetConfig.lookup.data.overallKeyDrivers.label
    description: @widgetConfig.lookup.data.overallKeyDrivers.description
    size: medium

    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }
    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.overallKeyDrivers.infoText
          label: @widgetConfig.lookup.data.overallKeyDrivers.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/score100"
      sortOrder: descending
      takeTop: 6
    }


   //filterexpression{ value: .dimension_score:dg1_dimensionScore = "Standard_3" }			

    row cut #itemsRow {
      total: none
      value: .item_score:dg1_questionScore
      //TODO: Need to exclude engagement items (filter out)
      // filter expression {
      //   value: .item_score:dg1_questionScore = "EV10137"      
      // }

    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:)
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint

        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }
    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }


    }



    column #gpr {
      label: "Percentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }


  widget dataGrid #overallTopPerform {
    label: @widgetConfig.lookup.data.overallTopPerform.label
    description: @widgetConfig.lookup.data.overallTopPerform.description
    size: medium
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.overallTopPerform.infoText
          label: @widgetConfig.lookup.data.overallTopPerform.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/gpr"
      sortOrder: descending
      takeTop: 5
    }




   //filterexpression{ value: .dimension_score:dg1_dimensionScore = "Standard_3" }			

    row cut #itemsRow {
      total: none
      value: .item_score:dg1_questionScore
      //TODO: Need to exclude engagement items (filter out)
      // filter expression {
      //   value: .item_score:dg1_questionScore = "EV10137"      
      // }

    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:)
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint
        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }

    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }


    }



    column #gpr {
      label: "Precentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }

  widget chart #keyDemoChartTop {
    label: "Top Performing Demographic Groups"// @widgetConfig.lookup.data.summaryMTVKeyDemo.label
    description: @widgetConfig.lookup.data.summaryMTVKeyDemo.description
    size: medium
    layout: vertical
    legend: bottomCenter

    axis category {
      textSize: 150

    }

    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }

    category cutByMulti {
      value: :keyDemoCalc
      sortBy: "/score"
      sortOrder: descending
      takeTop: 3
      //total: none

    }


    series #score {
      label: "Engagement mean score"
      value: IIF(count(:) > 5 AND count(:) / count(:, true, "__top") > 0.03, :dimensionScore())

    }

    axis primary #primaryAxis {
      maxValue: 5
      minValue: 0
      format: numberStatisticDefaultFormatter
    }
    axis secondary #secondaryAxis {
      hide: true
    }
  }

  widget chart #keyDemoChartBottom {
    label: "Bottom Performing Demographic Groups"//@widgetConfig.lookup.data.summaryMTVKeyDemo.label
    description: @widgetConfig.lookup.data.summaryMTVKeyDemo.description
    size: medium
    layout: vertical
    legend: bottomCenter
    axis category {
      textSize: 150
    }

    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }

    category cutByMulti {
      value: :keyDemoCalc
      sortBy: "/score"
      sortOrder: ascending
      takeTop: 3
      //total: none

    }


    series #score {
      label: "Engagement mean score"
      value: IIF(count(:) > 5 AND count(:) / count(:, true, "__top") > 0.03, :dimensionScore())


    }

    axis primary #primaryAxis {
      maxValue: 5
      minValue: 0
    }
    axis secondary #secondaryAxis {
      hide: true
    }
    removeEmptyCategories: true
  }


  widget dataGrid #overallAddDimensions {
    label: @widgetConfig.lookup.data.overallAddDimensions.label
    description: @widgetConfig.lookup.data.overallAddDimensions.description

    size: large
    filter expression {
      value: .dimensions:includeHXWidget
    }

    //Gets the overall data
    scope reportingHierarchy {
      reportingHierarchy: unitHierarchy
      nodes: AllData
    }

    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.overallAddDimensions.infoText
          label: @widgetConfig.lookup.data.overallAddDimensions.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }

    row list #dimensions {
      table: .dimensions:
      value: .dimensions:id
      total: none
    }

    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :dimensionScore()
        }
        statistic mean #sig {
          testingType: T
          argument: .dimension_score:dimensionScoreValue
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"
      }
    }

    column #main {
      label: "Mean score"
      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          //CNJ126 arrows ↑↓ or  ↑ ↓
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='font-size: 20px; color:{color};'>{arrow}</span>{asteric}</pre>"//To add Astric: 
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

        // tooltipFormatString: "<b style='font-size:20px'>{historyMean}</b><br>Historical Mean Score" + "<br><b style='font-size:20px'>{change}</b><br> vs " + @surveyToCompareWith.selectedLabel + "<br><span style='  height: 25px;  width: 25px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }
    column #benchmark {
      label: "Percentile"
      cell custom {
        lookup rank #rank {
          takeInArray: Per
          mode percentile {
          }
          source: benchmarks
          mapping header {
            header: dimensions
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :dimensionScore()
          formatter: rankFormatter
        }
        lookup value #mean {
          source: benchmarks
          mapping header {
            header: dimensions
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: mean
          formatter: scoreFormatter
        }
        formula #tooltip {
          value: IIF(score[column = /history.current] >= 0, "percentile rank in " + @defaultBenchmmark.selectedLabel + "<br>benchmark mean value " + mean[], "too few responses")
        }
        formatString: "{rank}"
        tooltipFormatString: "<span style='font-size:30px;'>{rank}</span><br>" + @defaultBenchmmark.selectedLabel + "<br><br><span style='font-size:20px;'>{mean}</span><br>" + @defaultBenchmmark.selectedLabel + " Mean Score "
      }
    }
    column #recoding {
      label: " "
      sortable: false
      cell custom {
        formatString: " "
      }
    }

  }
}

page #detailedSelectors {
  showPrintButton: false
  modal: true
  modalSize: large

  widget headline {
    container: container flex {
      area #all {
        display: flex
        flexDirection: column
        alignItems: "stretch"

        area #selectors {
          display: flex
          flexDirection: row
          justifyContent: "space-evenly"
          area #current {
            display: flex
            width: "30%"
            flexDirection: column
            alignSelf: "flex-start"
            alignItems: "flex-start"
            area #currentLabel {
            }
            area #currentColumns {
            }
          }
          area #history {
            display: flex
            width: "30%"
            flexDirection: column
            alignSelf: "flex-start"
            alignItems: "flex-start"
            area #historyLabel {
            }
            area #surveysList {
              height: 100px
              display: block
              overflow: auto
            }
            area #surveysColumns {
              borderTop: "double"
              paddingTop: 10px
            }
          }
          area #benchmarks {
            display: flex
            width: "30%"
            flexDirection: column
            alignSelf: "flex-start"
            alignItems: "flex-start"
            area #benchamrksLabel {
            }
            area #benchmarksList {
              height: 100px
              display: block
              overflow: auto
            }
            area #benchmarksColumns {
              borderTop: "double"
              paddingTop: 10px
            }
          }
        }
        area #buttons {
          display: flex
          flexDirection: row
          justifyContent: "flex-end"
          margin: 20px
        }
      }
    }
    tile text {
      areaId: currentLabel
      value: "Current results"
      style {
        fontWeight: "bold"
        fontSize: "larger"
      }
    }
    select #currentSurveySubColumns {
      areaId: currentColumns
      label: "Within current survey"
      mode: multi
      view list {
      }
      applyOnEvent: savedDetailedSelectors
      options: item {value: score label: 'Mean Score'},
      item {value: overall label: 'Overall Organization Score'},
      item {value: vsoverall label: 'vs. Overall Organization (difference)'},
      item {value: favorable label: 'Percent Favorable'},
      item {value: neutral label: 'Percent Neutral'},
      item {value: unfovarable label: 'Percent Unfovarable'},      
      item {value: distribution label: 'Response Distribution'},
      item {value: responses label: 'Responses'}
      defaultOption: @viewDefault.selected.current.defaultOption
      onDefaultChange: reset
    }

    tile text {
      areaId: historyLabel
      value: "History"
      style {
        fontWeight: "bold"
        fontSize: "larger"
      }
    }
    select #surveysList {
      areaId: surveysList
      mode: multi
      view list {
      }
      // view listBox {
      //   height: 200px
      //   column {
      //     label: "Surveys"
      //     value: "label"
      //   }
      // }
      applyOnEvent: savedDetailedSelectors
      options: @dtSurveys.forSelect.data
      defaultOption: @viewDefault.selected.history.defaultOption
      compareBy: this.trendOrder
      onDefaultChange: reset
    }
    select #surveyListSubColumns {
      areaId: surveysColumns
      mode: multi
      view list {
      }
      applyOnEvent: savedDetailedSelectors
      options: item {label: 'Mean Score' value: surveysScore },
      item {label: 'vs. History (difference)' value:surveysChange},
      item {label: 'vs. History (significance)' value: surveysSig},
      item {label: 'Overall Org Score' value: surveysOverall},
      item {label: 'Percent Favorable' value: surveysFavorable},
      item {label: 'Percent Neutral' value: surveysNeutral},
      item {label: 'Percent Unfavorable' value: surveysUnfovarable},
      item {label: 'Responses' value: surveysResponses}
      defaultOption: @viewDefault.selected.historySubColumns.defaultOption
      onDefaultChange: reset
    }

    tile text {
      areaId: benchamrksLabel
      value: "Benchmarks"
      style {
        fontWeight: "bold"
        fontSize: "larger"
      }
    }
    select #benchmarksList {
      areaId: benchmarksList
      mode: multi
      view list {
      }
      // view listBox {
      //   height: 251px
      //   column {
      //     label: "Benchmarks"
      //     value: "label"
      //   }
      // }
      applyOnEvent: savedDetailedSelectors
      options: @dtBenchmarks.forSelect.data
      defaultOption: @viewDefault.selected.benchmarks.defaultOption
      compareBy: this.idText
      onDefaultChange: reset
    }
    select #benchmarksListSubColumns {
      areaId: benchmarksColumns
      mode: multi
      view list {
      }
      applyOnEvent: savedDetailedSelectors
      options: item {label: 'Benchmark Mean Score' value: mean   },
      item {label: 'vs. Benchmark (Difference)' value: diff   },
      item {label: '10th Percentile' value: benchPercentile10},
      item {label: '25th Percentile' value: benchPercentile25},      
      item {label: '50th Percentile' value: benchPercentile50},
      item {label: '75th Percentile' value: benchPercentile75},
      item {label: '90th Percentile' value: benchPercentile90}
      defaultOption: @viewDefault.selected.benchmarkSubColumns.defaultOption
      onDefaultChange: reset
    }
    tile text {
      areaId: buttons
      value: "Apply and close"
      action sendEvent {
        name: 'savedDetailedSelectors'
      }
      action closeModal {
      }
      fontSize: 20
      style {
        paddingLeft: 20px
        paddingRight: 20px
        fontWeight: bold
        color: rgba(0, 0, 0, 0.664)
        textAlign: right
        backgroundColor: #ffffff
        borderStyle: solid
        borderColor: rgba(0, 0, 0, 0.664)
        borderWidth: thin
        borderRadius: 55px
      }
    }
  }
}

page #itemDetail {
  label: "Items"
  scope reportingHierarchy {
    reportingHierarchy: unitHierarchy
    mode: @rollupMode.selected.mode
  }


  widget headline #topSelectors {
    size: large

    container: container flex {
      display: flex
      flexDirection: row
      padding: 20px
      gap: 20px
      alignItems: center
    }

    select #rows {
      label: "Display"
      options: item { label:Nested value: both},
      item { label:Dimensions value:dimensions },
      item { label:Items value:items }
    }
    select #viewDefault {
      label: 'Select view'
      options: item {
        label: Standard 
        value: {
          current: {defaultOption: score, vsoverall, distribution, responses}
          history: {defaultOption: '2'}
          historySubColumns: {defaultOption: surveysScore}
          benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
          benchmarkSubColumns: {defaultOption: 'diff'}
        }
        code: default
      },
      item {
        label: 'Compare history' 
        value: {
          current: {defaultOption:  score, vsoverall, responses}
          history: {defaultOption: '2'}
          //history: {defaultOption: '2', '3', '4'} 
          //historySubColumns: {defaultOption: surveysScore, surveysChange, surveysSig}
          historySubColumns: {defaultOption: surveysScore, surveysFavorable}
          // benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
          // benchmarkSubColumns: {defaultOption: 'diff'}
          benchmarks: {defaultOption: 'none'}
          benchmarkSubColumns: {defaultOption: 'none'}
        }
        code: history
        },
      item {
        label: 'Compare Benchmarks' 
        value: {
          current: {defaultOption: distribution, score, vsoverall, responses}
          history: {defaultOption: '2'} 
          historySubColumns: {defaultOption: surveysScore, surveysFavorable}
          benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
          benchmarkSubColumns: {defaultOption: 'mean'}
        }
        code: benchmarks
      }
    }

    tile text #buttonTile {
      value: "More Options.."
      fontSize: 20
      navigateTo: detailedSelectors
      style {
        paddingLeft: 20px
        paddingRight: 20px
        fontWeight: bold
        color: rgba(0, 0, 0, 0.664)
        textAlign: right
        backgroundColor: #ffffff
        borderStyle: solid
        borderColor: rgba(0, 0, 0, 0.664)
        borderWidth: thin
        borderRadius: 55px
      }
    }
  }

  widget dataGrid #itemsDetailGrid {
    virtualize: true
    viaStrategy: shortest
    suppression recordsBase {
      threshold: @suppressionThreshold.selected
    }
    // filter expression {
	  //   value: left(.item_score:ev10039_path, 9) = "Overall->"
    // }
    // scope reportingHierarchy {
    //       reportingHierarchy: unitHierarchy
    //       nodes: AllData
    //     }
    // ignoreFilters: @switchDimensionsOrItems.selected
    // filter expression #dimensionIdFilter {
    //   value: IN(.dimensionItems:dimensionId, @sDims.selected)
    // }
    // filter expression #itemIdFilter {
    //   value: IN(.dimensionItems:questionId, @sItems.selected)
    // }

    // select #switchDimensionsOrItems {
    //   options: item {label: 'Filter by dimensions' value: itemIdFilter},
    //   item {label: 'Filter by items' value: dimensionIdFilter}
    // }
    // select #sItems {
    //   label: 'Items'
    //   options: @dtItems.forSelect.data
    //   mode: multi
    // }
    // select #sDims {
    //   label: 'Dimensions'
    //   options: @dtDimensions.forSelect2.data
    //   mode: multi
    // }
    size: large

    // select #rows {
    //   label: "Display"
    //   options: item { label:Nested value: both},
    //   item { label:Dimensions value:dimensions },
    //   item { label:Items value:items }
    // }

    // select #viewDefault {
    //   label: 'Select view'
    //   options: item {
    //     label: Default 
    //     value: {
    //       current: {defaultOption: score, vsOverall, distribution, responses}
    //       history: {defaultOption: '2'}
    //       historySubColumns: {defaultOption: surveysScore}
    //       benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
    //       benchmarkSubColumns: {defaultOption: 'diff'}
    //     }
    //     code: default
    //   },
    //   item {
    //     label: 'Compare history' 
    //     value: {
    //       current: {defaultOption:  score, vsOverall, responses}
    //       history: {defaultOption: '2'}
    //       //history: {defaultOption: '2', '3', '4'} 
    //       //historySubColumns: {defaultOption: surveysScore, surveysChange, surveysSig}
    //       historySubColumns: {defaultOption: surveysScore, surveysFavorable}
    //       // benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
    //       // benchmarkSubColumns: {defaultOption: 'diff'}
    //       benchmarks: {defaultOption: 'none'}
    //       benchmarkSubColumns: {defaultOption: 'none'}
    //     }
    //     code: history
    //     },
    //   item {
    //     label: 'Compare Benchmarks' 
    //     value: {
    //       current: {defaultOption: distribution, score, vsoverall, responses}
    //       history: {defaultOption: '2'} 
    //       historySubColumns: {defaultOption: surveysScore, surveysFavorable}
    //       benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
    //       benchmarkSubColumns: {defaultOption: 'mean'}
    //     }
    //     code: benchmarks
    //   }
    //   //,
    //   // item {
    //   //   label: 'Percentiles'
    //   //   value: {
    //   //     current: {defaultOption: distribution, score, vsoverall, responses}
    //   //     history: {defaultOption: '2'} 
    //   //     historySubColumns: {defaultOption: surveysScore}
    //   //     benchmarks: {defaultOption: @defaultBenchmmark.selected.idText  }
    //   //     benchmarkSubColumns: {defaultOption: 'benchPercentile10', benchPercentile50, benchPercentile75, benchPercentile90}
    //   //     }
    //   //     code: percentiles
    //   // }
    // }

    // select #currentSurveySubColumns {
    //   label: "Within current survey"
    //   mode: multi
    //   options: item {value: score label: 'Mean Score'},
    //   item {value: overall label: 'Overall Organization Score'},
    //   item {value: vsoverall label: 'vs. Overall Organization (difference)'},
    //   item {value: favorable label: 'Percent Favorable'},
    //   item {value: neutral label: 'Percent Neutral'},
    //   item {value: unfovarable label: 'Percent Unfovarable'},      
    //   item {value: distribution label: 'Response Distribution'},
    //   item {value: responses label: 'Responses'}
    //   defaultOption: @viewDefault.selected.current.defaultOption
    // }

    // select #surveysList {
    //   mode: multi
    //   label: "History"
    //   options: @dtSurveys.forSelect.data
    //   defaultOption: @viewDefault.selected.history.defaultOption
    //   compareBy: this.trendOrder
    // }
    // select #surveyListSubColumns {
    //   mode: multi
    //   label: 'Within history'
    //   options: item {label: 'Mean Score' value: surveysScore },
    //   item {label: 'vs. History (difference)' value:surveysChange},
    //   item {label: 'vs. History (significance)' value: surveysSig},
    //   item {label: 'Overall Org Score' value: surveysOverall},
    //   item {label: 'Percent Favorable' value: surveysFavorable},
    //   item {label: 'Percent Neutral' value: surveysNeutral},
    //   item {label: 'Percent Unfavorable' value: surveysUnfovarable},
    //   item {label: 'Responses' value: surveysResponses}
    //   defaultOption: @viewDefault.selected.historySubColumns.defaultOption
    // }
    // select #benchmarksList {
    //   mode: multi
    //   label: 'Benchmarks'
    //   options: @dtBenchmarks.forSelect.data
    //   defaultOption: @viewDefault.selected.benchmarks.defaultOption
    //   compareBy: this.idText
    // }
    // select #benchmarksListSubColumns {
    //   mode: multi
    //   label: 'Within benchmarks'
    //   options: item {label: 'Benchmark Mean Score' value: mean   },
    //   item {label: 'vs. Benchmark (Difference)' value: diff   },
    //   item {label: '10th Percentile' value: benchPercentile10},
    //   item {label: '25th Percentile' value: benchPercentile25},
    //   item {label: '50th Percentile' value: benchPercentile50},
    //   item {label: '75th Percentile' value: benchPercentile75},
    //   item {label: '90th Percentile' value: benchPercentile90}
    //   defaultOption: @viewDefault.selected.benchmarkSubColumns.defaultOption

    // }

    activeColumns: history, @currentSurveySubColumns.selected, surveys, bench
    activeRows: @rows.selected
    row nestedHeaders #both {
      viewMode: expanded
      nesting byTable {
        parent: .dimensionItems:dimensionId
        child: .dimensionItems:questionId
      }

      parent list #dimensions {
        total: none
        table: .dimensions:
        value: .dimensions:Id
        sortOrder: ascending
      }

      child list #items {
        total: none
        table: .items:
        value: toText(.items:SequenceId) + ".  " + answerText(.items:Id)
        sortBy: .items:SequenceId
        sortOrder: ascending
      }
    }
    row list #items {
      total: none
      table: .items:
      value: toText(.items:SequenceId) + ". " + answerText(.items:Id)
      sortBy: .items:SequenceId
      sortOrder: ascending
    }
    row list #dimensions {
      total: none
      table: .dimensions:
      value: .dimensions:Id
      sortOrder: ascending

    }

    column cutByTable #history {
      notAnswered: first

      //hide: true
      showLabel: true
      scope filter {
        name: period
        value: allDataHistory
      }
      total: none
      table: .reportHistory:

      column #historyMain {
        label: Main
      }
      column #historyOverall {

        label: Overall
        scope reportingHierarchy {
          reportingHierarchy: unitHierarchy
          nodes: AllData
        }
        scope filter {
          name: period
          value: allDataHistory
        }

        // filter expression {
        //   value: _isNotNull(@unitHierarchy.source)
        // }
      }
      column cut #historyDistributionDimensions {
        notAnswered: first
        total: none
        value: .dimension_score:threePoint
      }
      column cut #historyDistributionItems {
        notAnswered: first
        total: none
        value: .item_score:threePoint
      }
    }

    cell custom {
      row: dimensions
      column: historyOverall
      expression #score {
        value: :dimensionScore()
      }
      formatString: '{score}'
    }
    cell custom {
      row: items
      column: historyOverall
      expression #score {
        value: :itemScore() //:itemScoreSum() / :itemScoreCount()
      }
      formatString: '{score}'
    }

    cell custom {
      column: historyDistributionDimensions
      row: dimensions
      statistic percent #value {
        value: count(.dimension_score:)
        dimension: columns
      }
      formatString: "{value}"
    }
    cell custom {
      column: historyDistributionDimensions
      row: items
      formula #value {
        value: ''
      }
      formatString: '{value}'
    }
    cell custom {
      column: historyDistributionItems
      row: items
      statistic percent #value {
        value: count(.item_score:)
        dimension: columns
      }
      formatString: "{value}"
    }
    cell custom {
      column: historyDistributionItems
      row: dimensions
      formula #value {
        value: ''
      }
      formatString: '{value}'
    }
    column #overall {
      label: 'Overall'
    }
    column #distribution {
      label: "Response Distribution"
    }
    column #score {
      label: "Mean Score"
    }
    column #vsoverall {
      label: "vs Overall"
    }
    column #favorable {
      label: Favorable
    }
    column #neutral {
      label: Neutral
    }
    column #unfovarable {
      label: Unfovarable
    }

    cell custom {
      column: overall
      formula #score {
        value: score[column = /history.1/historyOverall]
        formatter: scoreFormatter
      }
      formatString: "{score}"
    }
    cell custom {
      column: vsoverall
      formula #vs {
        value: score[column = /history.1/historyMain] - score[column = /history.1/historyOverall]
        formatter: scoreFormatter
      }
      formatString: "{vs}"
    }
    //MG Need to hide if no previous survey but sould still be propeperly defined, May set previous as current
    // column #vsPrevious {
    //   label: "vs [default] " + @surveyToCompareWith.selectedLabel
    //   column #scorePrevious {
    //     label: "Mean score"
    //     cell custom {
    //       formula #score {
    //         value: score[column = /history.2/historyMain]
    //         formatter: floatDefaultFormatter
    //       }
    //       formatString: "{score}"
    //     }
    //   }
    //   column #diffPrevious {
    //     label: "Diff"
    //     cell custom {
    //       formula #diff {
    //         value: score[column = /history.1/historyMain] - score[column = /history.2/historyMain]
    //         formatter: floatDefaultFormatter
    //       }
    //       formatString: "{diff}"
    //     }
    //   }
    //   column #sigPrevious {
    //     label: "Sig"
    //     cell custom {
    //       formula #asteric {
    //         value: IIF(sig[column = /history.2/historyMain] != 0, "*", " ")
    //       }
    //       formatString: "{asteric}"
    //     }
    //   }
    // }

    cell microchart {
      row: items
      column: distribution
      value: count(.item_score:) + 3
      breakdownBy cut {
        value: .item_score:threePoint
      }
      microchart stacked100PercentBar {
        palette: favorable
      }
    }
    cell microchart {
      row: dimensions
      column: distribution
      value: count(.dimension_score:)  //count(:)
      breakdownBy cut {
        value: .dimension_score:threePoint
      }
      microchart stacked100PercentBar {
        palette: favorable
      }
    }
    cell custom {
      row: dimensions
      column: historyMain
      expression #score {
        value: :dimensionScore()
      }
      statistic mean #sig {
        testingType: T
        argument: .dimension_score:dimensionScoreValue
        compare: first
      }

      formula #diff {
        value: score[column = %.1] - score[]
      }
      formula #diffSum {
        value: sum(diff[column = %.*])
      }
      formula #count {
        value: count(score[column = %.*])
      }
      expression #responses {
        value: count(.dimension_score:)
      }
      formatString: "{score} [{sig}] {diffSum} {count} {responses}"

      tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}abc"
    }
    cell custom {

      row: items
      column: historyMain
      expression #score {
        value: :itemScore() // :itemScoreSum() / :itemScoreCount() // 
      }
      statistic mean #sig {

        testingType: T
        argument: numeric(.item_score:questionScoreValue)
        compare: first
      }

      formula #diff {
        value: score[column = %.current] - score[]
      }
      formula #diffSum {
        value: sum(diff[column = %.*])
      }
      formula #count {
        value: count(score[column = %.*])
      }
      expression #responses {
        value: count(.item_score:)
      }
      formatString: "{score} [{sig}] {diffSum} {count} {responses}"
      tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}abc"
    }
    cell custom {
      column: score
      formula #score {
        value: score[column = /history.1/historyMain]
        formatter: scoreFormatter
      }
      formatString: "{score}"
    }
    cell custom {
      column: favorable
      row: dimensions
      formula #value {
        value: value[column = /history.1/historyDistributionDimensions.1]
      }
      formatString: '{value}'
    }
    cell custom {
      column: neutral
      row: dimensions
      formula #value {
        value: value[column = /history.1/historyDistributionDimensions.2]
      }
      formatString: '{value}'
    }
    cell custom {
      column: unfovarable
      row: dimensions
      formula #value {
        value: value[column = /history.1/historyDistributionDimensions.3]
      }
      formatString: '{value}'
    }
    cell custom {
      column: favorable
      row: items
      formula #value {
        value: value[column = /history.1/historyDistributionItems.1]
      }
      formatString: '{value}'
    }
    cell custom {
      column: neutral
      row: items
      formula #value {
        value: value[column = /history.1/historyDistributionItems.2]
      }
      formatString: '{value}'
    }
    cell custom {
      column: unfovarable
      row: items
      formula #value {
        value: value[column = /history.1/historyDistributionItems.3]
      }
      formatString: '{value}'
    }




    column cutByTable #surveys {
      notAnswered: first
      scope filter {
        name: period
        value: AllPeriods
      }
      filter expression {
        value: IN(.reportHistory:historyTrendOrder, @surveysList.selected)
      }
      filter expression {
        value: .reportHistory:historyTrendOrder > 1

      }

      total: none
      table: .reportHistory:
      label: .reportHistory:historyLabel
      activeColumns: 'dummyInSurveys', @surveyListSubColumns.selected
      //MG have to include current as masking it out will totall exclude it from formulas
      //categories: "!'current'"
      column #dummyInSurveys {
        hide: true
        cell custom {
          formula #value {
            value: ''
          }
          formatString: ''
        }
      }
      column #surveysScore {
        label: "score"
        cell custom {
          formula #value {
            value: score[column = /history.%/historyMain]
          }
          formatString: '{value}'
        }
      }
      column #surveysChange {
        label: "change"
        cell custom {
          formula #value {
            value: score[column = /history.1/historyMain] - score[column = /history.%/historyMain]
          }
          formatString: '{value}'
        }
      }
      column #surveysSig {
        label: "sig"
        cell custom {
          formula #value {
            value: IIF(sig[column = /history.%/historyMain] != 0, "*", " ")
          }
          formatString: '{value}'
        }
      }
      column #surveysOverall {
        label: 'overall'
        cell custom {
          formula #value {
            value: score[column = /history.%/historyOverall]
          }
          formatString: '{value}'
        }
      }
      column #surveysResponses {
        label: 'responses'
        cell custom {
          formula #value {
            value: responses[column = /history.%/historyMain]
          }
          formatString: '{value}'
        }
      }
      column #surveysFavorable {
        label: Favorable
      }

      column #surveysNeutral {
        label: Neutral
      }

      column #surveysUnfovarable {
        label: Unfovarable
      }

    }
    cell custom {
      column: surveysFavorable
      row: dimensions
      formula #value {
        value: value[column = /history.%/historyDistributionDimensions.1]
      }
      formatString: '{value}'
    }
    cell custom {
      column: surveysNeutral
      row: dimensions
      formula #value {
        value: value[column = /history.%/historyDistributionDimensions.2]
      }
      formatString: '{value}'
    }
    cell custom {
      column: surveysUnfovarable
      row: dimensions
      formula #value {
        value: value[column = /history.%/historyDistributionDimensions.3]
      }
      formatString: '{value}'
    }
    cell custom {
      column: surveysFavorable
      row: items
      formula #value {
        value: value[column = /history.%/historyDistributionItems.1]
      }
      formatString: '{value}'
    }
    cell custom {
      column: surveysNeutral
      row: items
      formula #value {
        value: value[column = /history.%/historyDistributionItems.2]
      }
      formatString: '{value}'
    }
    cell custom {
      column: surveysUnfovarable
      row: items
      formula #value {
        value: value[column = /history.%/historyDistributionItems.3]
      }
      formatString: '{value}'
    }
    cell custom {
      row: items
      column: surveysScore
      expression #score {
        value: :itemScore() //:itemScoreSum() / :itemScoreCount() // :itemScore()
        formatter: scoreFormatter
      }

      formatString: "{score}"
    }
    cell custom {
      row: dimensions
      column: surveysScore
      expression #score {
        value: :dimensionScore()
        formatter: scoreFormatter
      }
      formatString: "{score}"
    }





    column cutByTable #bench {
      notAnswered: first
      table: .benchmarks:
      sortBy: .benchmarks:benchmarkOrder
      label: .benchmarks:benchmarkName
      filter expression {
        value: IN(.benchmarks:benchmarkID, @benchmarksList.selected)
      }
      activeColumns: 'dummyInBench', meanHidden, @benchmarksListSubColumns.selected
      column #dummyInBench {
        hide: true
        cell custom {
          formula #value {
            value: ''
          }
          formatString: ''
        }
      }
      column #meanHidden {
        label: "Mean hidden"
        hide: true
      }
      column #mean {
        label: "Mean"
      }
      column #diff {
        label: "Diff"
      }
      column #benchPercentile10 {
        label: '10th Percentile'
      }
      column #benchPercentile25 {
        label: '25th Percentile'
      }
      column #benchPercentile50 {
        label: '50th Percentile'
      }
      column #benchPercentile75 {
        label: '75th Percentile'
      }
      column #benchPercentile90 {
        label: '90th Percentile'
      }
    }
    cell custom {
      row: items
      column: benchPercentile90
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'items'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_90
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: dimensions
      column: benchPercentile90
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'dimensions'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_90
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: items
      column: benchPercentile75
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'items'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_75
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: dimensions
      column: benchPercentile75
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'dimensions'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_75
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: items
      column: benchPercentile25
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'items'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_25
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: dimensions
      column: benchPercentile25
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'dimensions'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_25
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: items
      column: benchPercentile50
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'items'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_50
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: dimensions
      column: benchPercentile50
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'dimensions'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_50
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: items
      column: benchPercentile10
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'items'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_10
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: dimensions
      column: benchPercentile10
      lookup value #value {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'dimensions'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Per_10
        formatter: scoreFormatter
      }
      formatString: '{value}'
    }
    cell custom {
      row: items
      column: meanHidden
      // expression #base {
      //   value: ""
      // }
      lookup value #mean {
        source: benchmarksById
        mapping header { //TODO: doesn't work yet, se comment on cutByTable #bench 
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'items'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Mean
        formatter: scoreFormatter
      }
      formatString: "{mean}"
    }
    cell custom {
      row: dimensions
      column: meanHidden
      // expression #base {
      //   value: ""
      // }
      lookup value #mean {
        source: benchmarksById
        mapping header {
          header: 'bench'
          selector: benchmarkID
        }
        mapping header {
          header: 'dimensions'
          selector: bmValueCode
        }
        // mapping value {
        //   selector: cmbdSurveyPID
        //   value: @externalConfig.combinedId
        // }
        value: Mean
        formatter: scoreFormatter
      }
      formatString: "{mean}"
    }
    cell custom {
      column: mean
      formula #mean {
        value: mean[column = /bench.%/meanHidden]
        formatter: scoreFormatter
      }
      formatString: "{mean}"
    }

    cell custom {
      column: diff
      formula #diff {
        value: score[column = /history.1/historyMain] - mean[column = /bench.%/meanHidden]
        formatter: scoreFormatter
      }
      formatString: "{diff}"
    }

    column #responses {
      label: "Responses"
      cell custom {
        expression #count {
          value: count(:)
        }
        formula #output {
          value: IIF(count[] < @suppressionThreshold.selected, "Too few responses", count[])
        }
        formatString: "{output}"
      }
    }


  }


}




page #orgDetails {
  label: "Work Units"
  scope reportingHierarchy {
    reportingHierarchy: unitHierarchy
    mode: @rollupMode.selected.mode
  }

  widget dataGrid {
    virtualize: true
    size: large
    select #rows {
      label: "Rows"
      options: item { label: "Nested mode" value: nested },
      item { label: "Flat mode" value: flat} 
    }
    select #sTMP {
      label: "Dimensions"
      mode: multi
      options: @dtDimensions.forSelect2.data
      defaultOption: true
      compareBy: this.isDefault
    }
    //MG might remove what is empty because of calculated value 
    //removeEmptyColumns: true
    filter expression {
      value: IN(.dimensions:id, @sTMP.selected)
    }
    suppression recordsBase {
      threshold: @suppressionThreshold.selected
    }
    activeRows: @rows.selected
    row comparison #nested {
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      reportingHierarchy: unitHierarchy
      mode: @rollupMode.selected.gridMode
      showTotal: true
      requestTotal: true
    }

    row comparisonFlat #flat {
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      reportingHierarchy: unitHierarchy
      labelStyle: nodeOnly
      showTotal: true
      mode: @rollupMode.selected.gridMode
    }
    column cutByTable #dimensions {
      table: .dimensions:
      hide: true
      scope filter {
        name: period
        value: allData
      }
      label: "to be hidden"
      showLabel: true
      total: none
      //value: .dimensions:id
      column cut #history {
        total: none
        value: .reportHistory:historyTypeCode
        cell custom {
          expression #score {
            value: :dimensionScore()
          }
          statistic mean #sig {
            testingType: T
            argument: .dimension_score:dimensionScoreValue
            compare: next
          }
          formula #diff {
            value: score[column = /dimensions.%/history.current] - score[]
            //MG this one shows strange results
            //value: score[column = /dimensions.%/history.current] - score[]
          }
          formula #diffSum {
            value: sum(diff[column = /dimensions.%/history.*])
          }
          formatString: "{score} [{sig}] {diff} {diffSum}"// {dummy}"
        }
      }
    }
    column cutByTable #engagement {
      showLabel: true
      table: .dimensions:
      //label: .dimensions:Label
      filter expression {
        value: .dimensions:isPrimary = true
      }
      column {
        label: "Mean Score"
        cell custom {
          formula #score {
            value: score[column = /dimensions.%/history.current]
          }
          formatString: "{score}"
        }
      }
      column {
        label: "Distribution"
        cell microchart {
          breakdownBy cut {
            value: .dimension_score:engagementFourPoint
          }
          value: :numberOfResponses()

          microchart stacked100PercentBar {
            palette: engaged
            //*NPL
            showLegend: true
          }
        }
      }
    }
    column cutByTable #team {
      showLabel: true
      table: .dimensions:
      //label: .dimensions:Label

      filter expression {
        value: .dimensions:id = "teamindex"
      }
      cell custom {
        formula #label {
          value: IIF(score[column = /dimensions.%/history.current] >= 4.15, "TI-1", IIF(score[column = /dimensions.%/history.current] < 3.80, "TI-3", IIF(score[column = /dimensions.%/history.current] > 3.80, "TI-2", "-")))
        }
        formatString: "{label}"
      }
    }

    column cutByTable #leader {
      showLabel: true
      table: .dimensions:
      //label: .dimensions:Label
      filter expression {
        value: .dimensions:id = "leaderindex"
      }
      cell custom {
        formula #label {
          value: IIF(score[column = /dimensions.%/history.current] >= 4, "High", IIF(score[column = /dimensions.%/history.current] <= 2.50, "Low", IIF(score[column = /dimensions.%/history.current] > 2.50, "Medium", "-")))
        }
        formatString: "{label}"
      }
    }
    column cutByTable #standard {
      showLabel: true
      table: .dimensions:
      //label: .dimensions:Label
      sortOrder: ascending
      //MG - sortBy below doesn't work
      //sortBy: .dimensions:Label
      filter expression {
        value: .dimensions:isPrimary = false AND _not(in(.dimensions:id, "leaderindex", "teamindex"))
      }
      cell custom {
        formula #change {
          value: diffSum[column = /dimensions.%/history.current]
          formatter: scoreFormatter
        }
        formula #arrow {
          //CNJ126 arrows ↑↓ or  ↑ ↓
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /dimensions.%/history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /dimensions.%/history.current] != 0, "change is statistically significant", "change is not statistically significant")
        }
        formula #score {
          value: score[column = /dimensions.%/history.current]
          formatter: scoreFormatter
        }
        //MG the next headerInfo -> Internal server Error
        headerInfo #rowCode {
          headerId: @rows.selected
          type: code
        }
        formula #vsOverall {
          value: IIF(rowCode[] != "__total__", score[] - score[row = %.__total__], " ")
          formatter: scoreFormatter
        }
        // formula #vsOverall {
        //   value: score[] - score[row = %.__total__]
        //   formatter: scoreFormatter
        // }
        formatString: "<pre>{score} {arrow}{asteric}<br>{vsOverall}   </pre>"
        tooltipFormatString: "change {change} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}" + "<br>vs Overall {vsOverall}"
      }
    }

    column #responses {
      label: "Responses"
      cell custom {
        expression #count {
          value: count(:)
        }
        formula #output {
          value: IIF(count[] < @suppressionThreshold.selected, "Too few responses", count[])
        }
        formatString: "{output}"
      }
    }
    column #isRollup {
      label: "Rollup"
      cell {
        value: IIF(_not(IsLeaf(unitHierarchy:^hierarchy)), "*")
      }
    }
  }



}
page #demographicDetails {
  label: "Demographics"
  scope reportingHierarchy {
    reportingHierarchy: unitHierarchy
    mode: @rollupMode.selected.mode
  }

  dataTable #dtDemoItems {
    dataGrid #dgDemoItems {

      filter expression {
        value: .demo_items:cmbdSurveyPID = @externalConfig.combinedId
      }

      //TODO: Only list demographics user have access to!
      row list #demos {
        total: none
        table: .demo_items:
        value: ""
        filter expression {
          //here should be filter end user specific
          value: .demo_items:demoPermissionTypeCode = "sensitive"
        }
      }
      column #main {
        cell custom {
          expression #id {
            value: .demo_items:itemID
          }
          expression #label {
            value: .demo_items:itemLabel
          }
          formatString: "{id} {label}"
        }
      }
    }
    map #forSelect {
      from: "demos"
      to: item {
        label: this.main.label
        value: this.main.id
      }
    }
  }

  widget dataGrid @externalConfig.demographicsRows {
    select #sDemos {
      mode: multi
      label: "select variables"
      options: @dtDemoItems.forSelect.data
    }
    activeRows: total, @sDemos.selected
    size: large
    row #total {
      label: "Grand Total"
    }


    column {
      label: "count"
      cell {
        value: count(:)
      }
    }
  }



}
page #commentAnalytics {
  label: "Comment Analytics"
  scope reportingHierarchy {
    reportingHierarchy: unitHierarchy
    mode: @rollupMode.selected.mode
  }



  widget headline #headlineWidget_4 {
      //label: "Select Open Ended Item"
    size: large
    select #questionSelect {
      label: "Select Open Ended Item"
      options: @dtOpenItems.forSelect.data
      mode: multi
    }
    tile text {
      value: " "
    }
  }

  filter expression {
    value: IN(textAnalyticsDataset.overallScore:variable, @questionSelect.selected)
  }

  widget headline #headlineWidget {
    dataSet: textAnalyticsDataset
    label: "Top Positive Topics"
    filter expression {
      value: :responseCategoryGroup() = "Positive"
    }

    tile grid #gridTile {
      row selectedFlat #topPositiveTopics_gridTile_row {
        reportingHierarchy: :categoryHierarchy
      }
      cell #topPositiveTopics_gridTile_column_cell {
        value: count(.analysisRecord:)
        format: bigNumberFormatter
      }
      column #topPositiveTopics_gridTile_column {
        hide: false
      }
      sort rows #topPositiveTopics_gridTile_sort {
        sortBy: "/topPositiveTopics_gridTile_column"
        sortOrder: "descending"
        takeTop: 5
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: hierarchy
        row: @topPositiveTopics_gridTile_row
        column: @topPositiveTopics_gridTile_column
        cell: @topPositiveTopics_gridTile_column_cell
        sort: @topPositiveTopics_gridTile_sort
      }
      tileStyle #tileStyle {
        bulletBackgroundColor: #34ae9a
        bulletTextColor: #ffffff
      }
    }
  }

  widget headline #topNegativeTopics {
    dataSet: textAnalyticsDataset
    label: "Top Negative Topics"
    filter expression {
      value: :responseCategoryGroup() = "Negative"
    }
    tile grid #gridTile {
      row selectedFlat #topNegativeTopics_gridTile_row {
        reportingHierarchy: :categoryHierarchy
      }
      cell #topNegativeTopics_gridTile_cell {
        value: :categoryResponseBase()
        format: bigNumberFormatter
      }
      column #topNegativeTopics_gridTile_column {
        hide: false
      }
      sort rows #topNegativeTopics_gridTile_sort {
        sortBy: "/topNegativeTopics_gridTile_column"
        sortOrder: "descending"
        takeTop: 5
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: hierarchy
        row: @topNegativeTopics_gridTile_row
        column: @topNegativeTopics_gridTile_column
        cell: @topNegativeTopics_gridTile_cell
        sort: @topNegativeTopics_gridTile_sort
      }
      tileStyle #tileStyle {
        bulletBackgroundColor: #d02625
        bulletTextColor: #ffffff
      }
    }
  }

  widget headline #topTopics {
    dataSet: textAnalyticsDataset
    label: "Top Topics"
    tile grid #gridTile {
      row selectedFlat #topTopics_gridTile_row {
        reportingHierarchy: :categoryHierarchy
      }
      cell #topTopics_gridTile_cell {
        value: :numberOfTaResponses()
        format: bigNumberFormatter
      }
      column #topTopics_gridTile_column {
        hide: false
      }
      sort rows #topTopics_gridTile_sort {
        sortBy: "/topTopics_gridTile_column"
        sortOrder: "descending"
        takeTop: 5
      }
      hint visualDesigner #visualDesignerHint {
        type: "rankedList"
        subType: hierarchy
        row: @topTopics_gridTile_row
        column: @topTopics_gridTile_column
        cell: @topTopics_gridTile_cell
        sort: @topTopics_gridTile_sort
      }
      tileStyle #tileStyle {
        bulletBackgroundColor: #576AD6
        bulletTextColor: #ffffff
      }
    }
  }


  widget hierarchyVisualization #hierarchyVisualizationWidget {
    dataSet: textAnalyticsDataset
    label: "Topic Hierarchy"
    size: large
    reportingHierarchy: textAnalyticsDataset:categoryHierarchy
    value size #sizeValue {
      value: textAnalyticsDataset:categoryResponseBase()
    }
    value color #colorValue {
      value: textAnalyticsDataset:categoryAverage()
      colorFormat: taSentimentColorFormatter
    }
    visualization treemap #treemapVisualization {
    }
  }

  widget dataGrid #dataGridWidget {
    dataSet: textAnalyticsDataset
    label: "Topic Explorer"
    size: large
    row comparison #comparisonRow {
      reportingHierarchy: :categoryHierarchy
    }

    column #copy_of_column_2 {
      label: "Percent of Total Responses"
      cell microchart #cell {
        format: percentDefaultFormatter
        value: :percentOfTaResponses()
        microchart bar #barMicrochart {
          max: 100
        }
      }
    }
    column #column_3 {
      label: "Number of Responses"
      cell #cell {
        value: :numberOfTaResponses()
        format: bigNumberFormatter
      }
    }
    column cut {
      value: :responseCategoryGroup()
      total: none

      cell columnPercentage #cell {
        value: :numberOfTaResponses()
      }
    }
    view comparativeStatistic #comparativeStatisticView {
      valueColorFormatter: taSentimentColorFormatter
      backgroundColorFormatter: taSentimentDefaultBackgroundColorFormatter
    }
    navigateTo: commentAnalyticsModal
  }
  config layout #layoutConfig {
    horizontalAlignmentMode: "threeColumnsCentered"
  }
}

page #comments {
  label: "Comments"
  hide: false
  modal: false

  widget comments #commentsWidget_3 {
    hide: true
    label: "Comments"
    column response #responseColumn {
      sortBy: comment
    }
    group question #questionGroup {
      label: "Comment"
      filter expression #excludeBlankResponses {
        value: :EV2023 != ""
      }
      comment: :EV2023
    }
    size: large
    table: :
    paginationType: paging
    showCountInLabel: true
    rowsPerPage: 50, 100, 200
  }

  widget comments #commentsWidget_2 {
    dataSet: textAnalyticsDataset
    label: "Comments"
    paginationType: paging
    showCountInLabel: true
    rowsPerPage: 50, 100, 200

    select #QuestionSelectCM {
      label: "Select open item"
      options: @dtOpenItems.forSelect.data
      mode: multi
    }

    overrideFilter level {
      name: "reportingHierarchyFilter"
      level: .overallScore:
      via: .categoryScore:
    }

    propagateFilter #propagateFilter {
      from: .model:
      to: .categoryScore:
      dropOriginal: true
    }
    propagateFilter #propagateFilter_2 {
      from: .categoryScore:
      to: .overallScore:
      dropOriginal: true
    }
    propagateFilter {
      from: .dimensionItems:
      to: .responseDimensions:
    }

    column response #responseColumn {
      sortBy: comment
      enableColumnFilter: false
    }
    group question #questionGroup {
      label: "Comment"
      filter expression #excludeBlankResponses {
        value: .overallScore:text != ""
      }
      comment: .overallScore:text
    }
    size: large
    table: .overallScore:
    navigateTo: TA_individualDetailsPage

    filter expression {
      value: IN(.overallScore:variable, @QuestionSelectCM.selected)

    }

    infobox #infobox {
      label: ""
      info: "Information here"
      size: "small"
    }
    cardAlign: none
  }

}


page #response_rates {

  widget chart #chartWidget {
    label: "Daily Response Count"
    animation: true
    series #series {
      chart area #barChart {
      }
      value: count(:responseid)
      format: bigNumberFormatter
      palette: defaultColorPalette
    }
    axis category #categoryAxis {
      axisLine: true
      tickLine: true
      textSize: 25
      orientation: -45
    }
    axis primary #primaryAxis {//hidden x
      hide: true
    }

    axis secondary #secondaryAxis { //hidden y
      hide: true

    }

    layout: "horizontal"
    size: large
    removeEmptyCategories: true

    category date #cutCategory {
      value: .response:interview_end
      breakdownBy: calendarDate
      format: dayformatter
    }

    series {
      label: ""
      value: parseInt("a")
      chart bar {
        legendType: none
      }
    }
    legend: "topLeft"
    description: "Tracking survey completions over time allows you to understand how many people on your team took time to complete the survey each day and are represented in the results."
    infobox #infobox {
      label: ""
      info: "Add text"
      size: "small"
    }
    cardShadow: false
  }


  widget dataGrid #dataGridWidget {
    virtualize: true
    select #rrRows {
      label: "Select Row"
      options: @dtResponseRateItems.forSelect2.data
    }
    activeRows: @rrRows.selected.row
    activeColumns: @rrRows.selected.col
    row comparison #hier {
      showTotal: false
      reportingHierarchy: unitHierarchy
    }
    row selectedFlat #units { //comparison {
      showTotal: false
      reportingHierarchy: unitHierarchy
      labelStyle: nodeOnly
    }
    row cut #cut {
      value: studio.expressionFromCdl(":" + @rrRows.selected.id)
    }

    column #invited {
      label: "Invited"
      cell {
        value: count(.respondent:, .respondent:Respondent = "Yes")
      }
    }
    column #responded {
      label: "Respondens"
      cell {
        value: count(:, :status = "complete")
      }
    }
    column #rate {
      label: "Response Rate"
      cell {
        value: formula {
          value: value[column = /responded] / value[column = /invited] * 100
        }
        format: percentDefaultFormatter
      }
    }
    column #rollup {
      label: "Rollup"
      cell {
        value: IIF(_NOT(isLeaf(unitHierarchy:^hierarchy)), "*")
      }
    }

    size: large
  }
  label: "Response Rates"
}


page #advanced_reporting {
  label: "Advanced Reporting"
  //replace with final version
  widget crosstab #crosstabWidget {
    size: "large"
    ignoreFilters: reportingPeriodFilter
    selectedSheet: "sheet_1"
    sheet #sheet_1 {
      name: "Sheet 1"
      scope reportingPeriod #reportingPeriodScope {
        period: AllData
      }
      settings #settings {
        nestSplits: true
        removeEmptyColumns: false
        columns splits #splitsColumns {
          column cut #cutColumn {
            value: :EV22642
            column cut #cutColumn_2 {
              value: :EV10020
              categories: "'1','2'"
              answersCount: 3
            }
            categories: "'1','2','3','4','5','6','7','8'"
            answersCount: 8
          }
        }
        rows questions #questionsRows {
          row cut #cutRow {
            value: :EV10234
          }
          row cut #cutRow_2 {
            value: :EV271
          }
        }
        transposed: false
        calculations #aC {
          calculation mean #meanCalculation {
            numberDecimals: 2
          }
          calculation categoricalMean #categoricalMeanCalculation {
            numberDecimals: 2
          }
        }
      }
      dataSet: surveyDataset
    }
  }
}

page #page_4 {
  hide: true
  label: "ConfigTest"
  widget markdown #markdownWidget {
    hide: @rolePermissions.permissionLookup.data.admin.isHidden
    label: "Needs admin permission"
    markdown: "Needs admin permission"
  }
  widget markdown #markdownWidget2 {
    hide: @rolePermissions.permissionLookup.data.summary.isHidden
    label: @widgetConfig.lookup.data.summaryMTVResponseRate.label
    description: @widgetConfig.lookup.data.summaryMTVResponseRate.description
    infobox {
      label: @widgetConfig.lookup.data.summaryMTVResponseRate.label
      info: @widgetConfig.lookup.data.summaryMTVResponseRate.infoText
    }
    markdown: "Widget needs summary permission"
  }
  widget dataGrid #dataGridWidget {
    label: "Permissions for role"
    size: "large"

    filter expression {
      value: .rolePermissions:cmbdSurveyPID = @externalConfig.combinedId AND .rolePermissions:roleCode = @userRole.selected
    }
    column #permissionCount {
      cell {
        value: count(.rolePermissions:permissionsCode)
      }
    }
    column #isHidden {
      label: "IsHidden"
      cell {
        value: count(.rolePermissions:permissionsCode) = 0
      }
    }
    row list #permissions {
      table: .allPermissions:
      value: .allPermissions:permissionsCode

    }


    //  map #forSelect {
    //   from: "permission"
    //   to: {
    //     permission: this.permission.value
    //   }
    // }
  }
  widget dataGrid #dataGridWidget_2 {
    label: "Data Grid"
    size: "large"
    filter expression {
      value: .rolePermissions:cmbdSurveyPID = @externalConfig.combinedId
    }
    column #widgetCode {
      cell {
        value: .widgetConfig:widgetCode
      }
    }
    column #widgetLabel {
      cell {
        value: .widgetConfig:widgetLabel
      }
    }
    column #widgetDescription {
      cell {
        value: .widgetConfig:widgetDescription
      }
    }
    column #widgetInfoText {
      cell {
        value: .widgetConfig:widgetInfoText
      }
    }
    row list #widgetCodes {
      table: .widgetConfig:
      value: .widgetConfig:widgetCode
    }
  }
  map #widgetConfigLookup {
    from: "widgetCodes"
    to:  {
      label: this.widgetLabel.value
      descripton: this.widgetDescription.value
      infoText: this.widgetInfoText.value
    }
    toRecord byKey {
      key: this.widgetCode.value
    }
  }
  widget table #tableWidget {
    label: "Dimensions"
    size: "large"
    table: .dimension_group_dimensions:
    showCodeLabelSelector: true
    column value #valueColumn {
      label: "id"
      value: .dimension_group_dimensions:id
      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "type"
      value: .dimension_group_dimensions:type
      enableColumnFilter: true
    }
  }

  widget dataGrid #dgDimensions {
    size: large
    row list #dimensions {
      total: none
      table: .dimensions:
      value: ""
      sortBy: "/_label"
      sortOrder: ascending
    }
    column #_label {
      hide: true
      cell {
        value: .dimensions:id //concatinate to force id instead of label
      }
    }
    column #results {
      cell custom {
        formula #label {
          value: [column = /_label]
        }
        expression #type {
          value: "leader" //.dimensions:typeMG
        }
        expression #id {
          value: toText(.dimensions:id)
        }
        expression #isDefault {
          value: .dimensions:isPrimary
        }
        formula #points {
          value: IIF(type[] = "Engagement", "fourPoint", "threePoint")
        }
        formatString: "{id}"
          //formatString: "{label} | {type} | {id} | {isDefault}"
      }
    }
  }
}
page #page_6 {
  hide: true
  label: "Page 6"

  widget dataGrid {
    label: "Item details"
    virtualize: true
    suppression recordsBase {
      threshold: @suppressionThreshold.selected
    }
    size: large
    select #rows {
      options: item { label:Nested value: both},
      item { label:Dimensions value:dimensions },
      item { label:Items value:items }
    }
    activeRows: @rows.selected

    row nestedHeaders #both {
      viewMode: expanded
      nesting byTable {
        parent: .dimensionItems:dimensionId
        child: .dimensionItems:questionId
      }

      parent list #dimensions {
        total: none
        table: .dimensions:
        value: .dimensions:Id
        sortOrder: ascending
      }

      child list #items {
        total: none
        table: .items:
        value: toText(.items:SequenceId) + ". " + answerText(.items:Id)
        sortBy: .items:SequenceId
        sortOrder: ascending
      }
    }
    row list #items {
      total: none
      table: .items:
      value: toText(.items:SequenceId) + ". " + answerText(.items:Id)
      sortBy: .items:SequenceId
      sortOrder: ascending
    }
    row list #dimensions {
      total: none
      table: .dimensions:
      value: .dimensions:Id
      sortOrder: ascending
    }

    // row #items {
    // }
    // row #dimensions {
    // }
    column cut #history {
      label: "Will be hidden"
      showLabel: true
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
    }
    column #overall {
      hide: true
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
    }
    column #distribution {
      label: "Response Distribution"
    }


    cell microchart {
      row: items
      column: distribution
      value: count(:) + 1
      breakdownBy cut {
        value: .item_score:threePoint
      }
      microchart stacked100PercentBar {
        palette: favorable
      }
    }



  }

  widget dataGrid #dgEngagementSummary {
    size: large
    filter expression {
      value: _isNotNull(@unitHierarchy.source)
    }
    suppression recordsBase {
      threshold: @suppressionThreshold.selected
    }

    row #engagement {
      filter expression {
        value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
      }
    }

    column cut #history {
      scope filter {
        name: period
        value: currentAndPrevious
      }
      value: .reportHistory:historyTypeCode
      total: none

      cell custom {
        expression #score {
          value: :dimensionScore()
            //formatter: numberFormatter_5
        }
        statistic mean #sig {
          testingType: T
          argument: .dimension_score:dimensionScoreValue
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diff}"
      }
    }
    column #main {
      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
        }
        formula #sig {
          value: sig[column = /history.current]
        }
        formula #asteric {
          value: IIF(sig[] != 0, "*", " ")
        }
        formula #arrow {
          //CNJ126 arrows ↑↓ or  ↑ ↓
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #sigInfo {
          value: IIF(sig[] != 0, "change is statistically significant", "change is not statistically significant")
        }
        formatString: "{current} ({change}) [{sig}]"
      }
    }

    column #benchmark {
      cell custom {
        lookup rank #rank {
          takeInArray: Per
          mode percentile {
          }
          source: benchmarks
          mapping value {
            value: @externalConfig.primaryDimensionId
            selector: bmValueCode
          }
            // mapping value { //TODO: 
            //   value: @defaultBenchmmark.selected.definitionId
            //   selector: DefinitionId
            // }
            // mapping value { //TODO: need trendYear in benchmark_values
            //   value: @defaultBenchmmark.selected.periodId
            //   selector: Period
            // }
          value: :dimensionScore()
          formatter: rankFormatter
        }
        formatString: "{rank}"
      }
    }
    column #microchart {
      cell microchart {
        value: count(.dimension_score:)
        breakdownBy cut {
          value: .dimension_score:engagementFourPoint
        }
        microchart pie {
        }
      }
    }
  }


  widget table #tableWidget {
    label: "Table"
    size: "large"
    table: .dimension_group_dimensions:
    showCodeLabelSelector: true
    column value #valueColumn {
      label: "description"
      value: .dimension_group_dimensions:description
      enableColumnFilter: true
    }
    column value #valueColumn_2 {
      label: "id"
      value: .dimension_group_dimensions:id
      enableColumnFilter: true
    }
    column value #valueColumn_3 {
      label: "includeHXWidget"
      value: .dimension_group_dimensions:includeHXWidget
      enableColumnFilter: true
    }
    column value #valueColumn_4 {
      label: "isPrimary"
      value: .dimension_group_dimensions:isPrimary
      enableColumnFilter: true
    }
    column value #valueColumn_5 {
      label: "parentDimension"
      value: .dimension_group_dimensions:parentDimension
      enableColumnFilter: true
    }
    column value #valueColumn_6 {
      label: "sequenceId"
      value: .dimension_group_dimensions:sequenceId
      enableColumnFilter: true
    }
    column value #valueColumn_7 {
      label: "type"
      value: .dimension_group_dimensions:type
      enableColumnFilter: true
    }
  }
  widget dataGrid #dgDimensions {
    size: large
    row list #dimensions {
      total: none
      table: .dimensions:
      value: ""
      sortBy: "/_label"
      sortOrder: ascending
    }
    column #_label {
        //hide: true
      cell {
        value: .dimensions:id
      }
    }
    column #results {
      cell custom {
        formula #label {
          value: [column = /_label]
        }
        expression #type {
          value: .dimensions:id //"leader" //.dimensions:typeMG
        }
        expression #id {
          value: .dimensions:id
        }
        expression #isDefault {
          value: .dimensions:isPrimary
        }
        formula #points {
          value: IIF(type[] = "Engagement", "fourPoint", "threePoint")
        }
        formatString: "{label} | {type} | {id} | {isDefault}"
      }
    }
  }
  widget table #tableWidget_2 {
    label: "Table"
    size: "large"
    table: .dg1_dimensionScore:
    column value #valueColumn {
      label: "combined_sourceid"
      value: .dg1_dimensionScore:combined_sourceid
      enableColumnFilter: true
    }
    column value #valueColumn {
      label: "combined_sourceid"
      value: .dg1_dimensionScore:reportHistoryId
      enableColumnFilter: true
    }
    column value #valueColumn2 {
      label: "ev10039"
      value: .dg1_dimensionScore:ev10039
      enableColumnFilter: true
    }
  }
}
page #page_12 {
  hide: true
  label: "Issues"
  widget chart #summaryMTVTrend {
    label: @widgetConfig.lookup.data.summaryMTVTrend.label
    description: @widgetConfig.lookup.data.summaryMTVTrend.description
    hide: @rollupMode.selected.mode != "rollup"

    scope filter {
      name: period
      value: AllPeriods
    }

    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }

    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVTrend.infoText
          label: @widgetConfig.lookup.data.summaryMTVTrend.label
        }
      }
      button #export {
        action export {
          format: png
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }

      // filter expression {
      //   value: .periods:includeInTrend
      // }
    filter expression {
      value: .dimension_score:dg1_dimensionScore = @externalConfig.primaryDimensionId
    }
    category cut #periods {
      value: .reportHistory:trendYear
      sortBy: .reportHistory:trendYear
      sortOrder: ascending
    }

    series {
      label: ""
      value: parseInt("a")
      chart bar {
        legendType: none
      }
    }
    // category list #periods {
    //   value: .reportHistory:historyLabel
    //   table: .reportHistory:
    //   sortBy: .reportHistory:historyTrendOrder

    //   sortOrder: ascending //TODO: sorting does not seem to work
    // }

    axis category {
      interval: preserveStartEnd
    }

    series #user {
      label: @rollupMode.selectedLabel
      value: :dimensionScore()
      chart line {
      }
    }
    series #entire {
      label: "Entire Organization"
      scope reportingHierarchy {
        reportingHierarchy: unitHierarchy
        nodes: AllData
      }
      filter expression {
        value: _isNotNull(@unitHierarchy.source)
      }
      value: :dimensionScore()
      chart line {
      }
    }
    series #benchm {

      label: @defaultBenchmmark.selected.definitionName
      value: lookup value {
        source: benchmarks
        mapping value {
          value: @externalConfig.primaryDimensionId
          selector: bmValueCode
        }
        mapping value {
          value: @defaultBenchmmark.selected.definitionId
          selector: benchmarkDefinitionID
        }
        mapping header {
          header: periods
          //value: .reportHistory:trendYear
          selector: TrendYear
        }
        value: mean
        formatter: scoreFormatter
      }
      chart line {
      }
    }
    legend: bottomCenter
    axis primary {
    }

    size: large
    axis secondary #secondaryAxis {
      hide: true
    }
  }
}
page #commentAnalyticsModal {
  // label: "Page 12"
  hide: false
  modal: true
  widget comments #comments3 {
    exportable: true
    table: textAnalyticsDataset.overallScore:
    label: "Comments"
    size: large
    showHeader: true
    sortOrder: ascending
    sortColumn: comments
    headerNumberOfLines: 3
    // navigateTo: Response
    stretchColumns: true
    paginationType: paging
    rowsPerPage: 100,150,250,500


    view metric #sentimentperformance {
      valueColorFormatter: sentimentindicatortext
      fontSize: small
      backgroundColorFormatter: sentimentindicator
    }
    view comment #viewComments {
      lines: 10
    }

    column response #comments {
      footer: surveyDataset.response:interview_start
      //header: @FieldsExit.CommentHeaderText
      view: viewComments
      width: 1000px
      enableColumnFilter: true
    }

    group question {
      label: "All Comments"
      comment: textAnalyticsDataset.overallScore:text

      column value {
        value: textAnalyticsDataset.overallScore:variable
        label: "Comment Field"
        enableColumnFilter: true
        width: 250px
        align: center
      }
      column metric #overallSentiment {
        label: "Overall Sentiment"
        value: textAnalyticsDataset:overallAverage()
        format: sentimentindicatortextValue
        target: 1
        view: sentimentperformance
        width: 120px
        align: center

      }
    }
    filter expression {
      value: surveyDataset:EV10040 != "" AND surveyDataset:respondent = "Yes" AND IN(textAnalyticsDataset.overallScore:variable, @questionSelect.selected)

    }

  }
}

page #page_16 {
  label: "Page 16"
  widget dataGrid #summaryMTVKeyDrivers {
    label: @widgetConfig.lookup.data.summaryMTVKeyDrivers.label
    description: @widgetConfig.lookup.data.summaryMTVKeyDrivers.description
    size: large
    hide: @rollupMode.selected.mode != "rollup"
    suppressRule {
      criteria: count(:, .reportHistory:historyTypeCode = "current") < 29999 + @suppressionThreshold.selected //when
      label: "The number of responses for your team is below the minimum threshold required to display results." //what to display
    }


    primaryBenchmarkId: @defaultBenchmmark.selected.idInt
    toolbar { // This 
      button #infobox {
        action showInfobox {
          size: large
          info: @widgetConfig.lookup.data.summaryMTVKeyDrivers.infoText
          label: @widgetConfig.lookup.data.summaryMTVKeyDrivers.label
        }
      }
      button #export {
        action export {
          format: default
        }
      }

      button #navigate {

        action navigate {
          navigateTo: itemDetails
        }

      }
    }
    filter expression {
      value: _isNotNull(:forDimension)

    }

    sort rows {
      sortBy: "/score100"
      sortOrder: descending
      takeTop: 6
    }


   //filterexpression{ value: .dimension_score:dg1_dimensionScore = "Standard_3" }			
    filter expression {
      value: .scaled_items:includeKD
    }

    row cutByTable #itemsRow {
      total: none
      table: .items:
    }

    column {
      label: "Response Distribution"
      cell microchart {
        row: items
        column: distribution
        value: count(:) + 1
        format: bigNumberFormatter
        breakdownBy cut {
          value: .item_score:threePoint

        }
        microchart stacked100PercentBar {
          palette: favorable


        }
      }
    }
    column cut #history {
      hide: true
      scope filter {
        name: period
        value: currentAndPrevious
      }
      total: none
      value: .reportHistory:historyTypeCode
      cell custom {
        expression #score {
          value: :itemScore()
        }
        statistic mean #sig {
          testingType: T
          argument: numeric(.item_score:questionScoreValue)
          compare: next
        }
        formula #diff {
          value: score[column = %.current] - score[]
        }
        formula #diffSum {
          value: sum(diff[column = %.*])
        }
        formatString: "{score} [{sig}] {diffSum}"
        tooltipFormatString: "{diff} vs " + @surveyToCompareWith.selectedLabel + "<br>{sigText}"

      }
    }
    column #main {
      label: "Mean Score"


      cell custom {
        formula #current {
          value: score[column = /history.current]
        }
        formula #change {
          value: diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }
        formula #arrow {
          value: IIF(change[] > 0, "↑", IIF(change[] < 0, "↓", "-"))
        }
        formula #asteric {
          value: IIF(sig[column = /history.current] != 0, "*", " ")
        }
        formula #sigText {
          value: IIF(sig[column = /history.current] != 0, "The change is statistically significant", "The change is not statistically significant")
        }
        formula #color {
          value: IIF(change[] > 0, IIF(sig[column = /history.current] != 0, "#34ae9a", "Black"), IIF(change[] < 0, IIF(sig[column = /history.current] != 0, "#d02625", "Black"), "Black"))
        }
        formula #historyMean {
          value: score[column = /history.current] - diffSum[column = /history.current]
          formatter: floatDefaultFormatter
        }

        formatString: "<pre>{current}<span style='color:{color};font-size:20px'>{arrow}</span>{asteric}</pre>"
        tooltipFormatString: "<span style='font-size:30px'>{historyMean}</span><br>Historical Mean Score" + "<br><br><span style='font-size:20px'>{change}</span><br> vs " + @surveyToCompareWith.selectedLabel + "<br><br><span style='  height: 15px;  width: 15px;  background-color: {color};  border-radius: 50%;  display: inline-block;' class='dot'></span><br>{sigText}"

      }
    }

    //column cut {value: .dimension_score:dg1_dimensionScore }
    column #cof {
      hide: true
      label: "Correlation"
      cell {
        value: correlation(score(.item_score:questionScoreValue), :forDimension)
      }
    }
    column #corHundred {
      hide: true
      label: "Correlation Scale100"
      cell custom {
        //ScaledValue = (v - MIN(AllValues)) / (MAX(AllValues) - MIN(AllValues)) * (SCALE_MAX - SCALE_MIN) + SCALE_MIN
        formula #max {
          value: max(value[row = /itemsRow.*, column = /cof])
        }
        formula #min {
          value: min(value[row = /itemsRow.*, column = /cof])
        }
        formula #coefficient {
          value: value[column = /cof]
        }
        formula #scaled100 {
          value: (coefficient[] - min[]) / (max[] - min[]) * 100
        }

        formatString: "{scaled100}"
      }


    }



    column #gpr {
      label: "Percentile"
      cell {
        value: lookup rank {
          takeInArray: Per

          mode percentile {

          }
          source: benchmarks
          mapping header {
            header: itemsRow
            selector: bmValueCode
          }
          mapping value {
            value: @defaultBenchmmark.selected.definitionId
            selector: BenchmarkDefinitionId
          }

          mapping value {
            value: @defaultBenchmmark.selected.periodId
            selector: TrendYear
          }
          value: :itemScore()
        }
        format: rankFormatter

      }

    }
    column #addtoPlan {
    // hide: true
      label: "Add to Plan"
      cell {
        value: "+"

      }

    }

    column #score100 {
      hide: true
      label: "Score100"
      cell {
        value: formula {
          value: scaled100[column = /corHundred] - value[column = /gpr]
        }

      }
    }
  }
}
